

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
Use ieee.std_logic_arith.all;
Use ieee.std_logic_unsigned.all;


entity MUX_signal_type_PP is

	generic (
	
	  data_pft: integer := 6;
		data_ppz : integer := 5;
		data_rom : integer := 14
				);
	Port(
		Clk_96 : in std_logic;
		Ce_F6 : in std_logic;
		En : in std_logic;
		OD : in std_logic;		
	   LG : in std_logic;		
	   TI : in std_logic;
		fdop	  : in std_logic_vector (7 downto 0);
		fdev	: in std_logic_vector (2 downto 0);  
		ppz_m : in std_logic_vector (4 downto 0);
		PFT : in std_logic_vector (data_pft downto 1);
		pipp : in std_logic;
		--P2 : in std_logic_vector (1 downto 0);

		--NT_PPZ : in std_logic_vector (data_ppz downto 1);----------?
		Sign_LCHM : in std_logic;

		Rom_cos : out std_logic_vector (data_rom-1 downto 0)
		--Rom_cos : out std_logic_vector (7 downto 0)
	);

end MUX_signal_type_PP;

architecture Behavioral of MUX_signal_type_PP is

--Signal P1_P2_PFT : std_logic_vector(5 downto 1):=(others => '0');
	signal P2_PFT : std_logic_vector(data_pft downto 1):=(others => '0');
	
	signal Rom_cos_L7C3_i : integer;
	signal Rom_cos_L7C4_i : integer;
	signal Rom_cos_L11C3_i : integer;
	signal Rom_cos_L11C4_i : integer;
	signal Rom_cos_L15C3_i : integer;
   signal Rom_cos_L15C4_i : integer;
   signal Rom_cos_L19C3_i : integer;
	signal Rom_cos_L23C3_i : integer;
   signal Rom_cos_L23C4_i : integer;
	signal Rom_cos_L11_i : integer;
	signal Rom_cos_L15_i : integer;
	signal Rom_cos_L23_i : integer;
	signal Rom_cos_L30_i : integer;
	signal Rom_cos_L3_plus : integer;
	signal Rom_cos_L3_minus : integer;

  signal Rom_cos_out : std_logic_vector (data_rom-1 downto 0):=(others => '0');
--Signal Rom_sin_i : integer range -64 to 64;
--Signal Rom_cos_i : integer range -64 to 64;
	signal Rom_cos_i : integer;

begin



--------------------------------  L ������ '+'
LHM_PP2: entity work.LHM_ALL
generic map(

		rom_cos =>
		--(100, 8185, 702, -8117, -1499, 7969, 2280, -7746, -3040, 7447, 3770, -7079, -4464, 6640, 5114, -6140, -5716, 5580, 6262, -4967, -6749, 4306, 7170, -3605, -7523, 2868, 7803, -2105, -8010, 1321, 
--8138, -526, -8191, -275, 8163, 1072, -8059, -1860, 7876, 2629, -7620, -3374, 7290, 4085, -6892, -4758, 6427, 5384, -5903, -5961, 5320, 6479, -4689, -6937, 4012, 7328, -3299, -7650, 2552, 7898, 
---1784, -8072, 996, 8169, -202, -8189, -596, 8130, 1387, -7996, -2166, 7784, 2922, -7501, -3653, 7145, 4346, -6723, -5001, 6236, 5606, -5693, -6160, 5093, 6654, -4448, -7087, 3759, 7451, -3036, 
---7746, 2284, 7967, -1512, -8115, 723, 8184, 69, -8178, -863, 8094, 1647, -7935, -2417, 7700, 3162, -7394, -3879, 7018, 4558, -6578, -5195, 6074, 5782, -5515, -6317, 4903, 6790, -4247, -7202, 
--3550, 7544, -2821, -7818, 2065, 8016, -1291, -8142, 503, 8190, 287, -8163, -1076, 8058, 1853, -7880, -2614, 7627, 3349, -7305, -4055, 6913, 4721, -6459, -5344, 5942, 5916, -5373, -6435, 4752, 
--6892, -4089, -7287, 3386, 7612, -2654, -7868, 1896, 8050, -1122, -8159, 336, 8190, 450, -8148, -1235, 8028, 2006, -7836, -2760, 7570, 3486, -7236, -4183, 6833, 4838, -6370, -5451, 5846, 6011, 
---5270, -6517, 4643, 6962, -3976, -7344, 3271, 7657, -2538, -7901, 1779, 8071, -1007, -8168, 223, 8189, 560, -8136, -1341, 8007, 2106, -7806, -2854, 7532, 3574, -7191, -4263, 6782, 4911, -6313, 
---5516, 5785, 6068, -5206, -6566, 4578, 7003, -3910, -7377, 3204, 7682, -2471, -7919, 1714, 8082, -944, -8173, 163, 8187, 617, -8129, -1393, 7996, 2155, -7791, -2898, 7514, 3613, -7171, -4297, 
--6760, 4940, -6291, -5540, 5762, 6088, -5184, -6582, 4556, 7015, -3890, -7386, 3186, 7688, -2456, -7923, 1702, 8083, -935, -8173, 157, 8187, 620, -8129, -1393, 7996, 2151, -7793, -2892, 7517, 
--3604, -7176, -4286, 6769, 4927, -6302, -5526, 5778, 6073, -5203, -6567, 4580, 7000, -3917, -7372, 3218, 7676, -2492, -7913, 1742, 8076, -979, -8170, 205, 8188, 569, -8136, -1340, 8008, 2096, 
---7811, -2835, 7542, 3547, -7208, -4229, 6807, 4871, -6348, -5471, 5831, 6021, -5263, -6519, 4647, 6956, -3992, -7334, 3299, 7644, -2579, -7888, 1834, 8060, -1076, -8162, 306, 8190, 465, -8147, 
---1233, 8030, 1988, -7844, -2728, 7586, 3441, -7263, -4125, 6874, 4771, -6427, -5376, 5920, 5932, -5364, -6437, 4758, 6883, -4112, -7270, 3428, 7591, -2716, -7847, 1979, 8032, -1226, -8148, 460, 
--8190, 307, -8162, -1074, 8061, 1828, -7890, -2569, 7649, 3285, -7342, -3974, 6968, 4625, -6536, -5238, 6045, 5803, -5503, -6319, 4910, 6778, -4277, -7179, 3605, 7515, -2903, -7787, 2174, 7990, 
---1428, -8124, 668, 8185, 95, -8178, -860, 8096, 1615, -7946, -2358, 7725, 3078, -7439, -3773, 7086, 4433, -6674, -5056, 6202, 5633, -5678, -6163, 5102, 6638, -4485, -7056, 3827, 7412, -3138, 
---7705, 2419, 7929, -1682, -8087, 929, 8172, -170, -8189, -593, 8133, 1348, -8008, -2093, 7813, 2818, -7552, -3520, 7224, 4190, -6836, -4826, 6387, 5418, -5885, -5965, 5331, 6459, -4732, -6899, 
--4092, 7277, -3418, -7595, 2713, 7845, -1987, -8030, 1242, 8145, -489, -8191, -271, 8165, 1026, -8071, -1773, 7906, 2504, -7675, -3215, 7377, 3896, -7017, -4546, 6596, 5155, -6121, -5721, 5591, 
--6237, -5016, -6701, 4397, 7106, -3741, -7452, 3053, 7733, -2340, -7950, 1606, 8097, -860, -8177, 105, 8186, 648, -8127, -1398, 7997, 2134, -7802, -2854, 7538, 3547, -7212, -4212, 6824, 4839, 
---6380, -5427, 5879, 5966, -5332, -6458, 4737, 6892, -4104, -7270, 3435, 7585, -2739, -7838, 2018, 8022, -1283, -8141, 534, 8189, 216, -8170, -967, 8080, 1707, -7925, -2435, 7701, 3140, -7414, 
---3820, 7063, 4467, -6654, -5077, 6188, 5643, -5673, -6163, 5107, 6630, -4502, -7043, 3856, 7395, -3181, -7686, 2477, 7912, -1754, -8073, 1015, 8165, -270, -8191, -479, 8146, 1222, -8035, -1957, 
--7856, 2673, -7613, -3369, 7305, 4034, -6937, -4668, 6511, 5261, -6032, -5812, 5501, 6312, -4927, -6762, 4310, 7154, -3660, -7488, 2977, 7758, -2272, -7966, 1546, 8105, -809, -8180, 64, 8185, 
--679, -8124, -1419, 7994, 2144, -7800, -2854, 7540, 3538, -7219, -4195, 6838, 4815, -6401, -5397, 5911, 5932, -5373, -6420, 4790, 6854, -4170, -7233, 3513, 7550, -2829, -7808, 2121, 7999, -1397, 
---8126, 660, 8185, 80, -8179, -821, 8104, 1553, -7964, -2275, 7758, 2976, -7489, -3654, 7158, 4300, -6770, -4913, 6326, 5483, -5831, -6011, 5287, 6487, -4703, -6913, 4078, 7280, -3422, -7590, 
--2736, 7835, -2030, -8019, 1306, 8136, -574, -8189, -165, 8173, 901, -8093, -1630, 7945, 2345, -7735, -3042, 7460, 3713, -7127, -4355, 6734, 4960, -6289, -5526, 5791, 6046, -5249, -6519, 4662, 
--6937, -4040, -7300, 3383, 7603, -2701, -7847, 1996, 8025, -1277, -8141, 545, 8189, 188, -8173, -922, 8089, 1646, -7942, -2359, 7730, 3051, -7458, -3720, 7124, 4357, -6734, -4961, 6289, 5523, 
---5796, -6042, 5254, 6511, -4673, -6930, 4052, 7292, -3401, -7597, 2722, 7839, -2022, -8020, 1305, 8136, -579, -8189, -153, 8174, 882, -8096, -1605, 7952, 2313, -7747, -3005, 7478, 3671, -7152, 
---4309, 6767, 4911, -6330, -5476, 5841, 5996, -5308, -6469, 4731, 6889, -4119, -7257, 3472, 7565, -2801, -7815, 2105, 8001, -1394, -8126, 671, 8185, 55, -8181, -783, 8110, 1502, -7978, -2212, 
--7780, 2901, -7524, -3570, 7206, 4208, -6834, -4815, 6406, 5382, -5930, -5909, 5405, 6387, -4840, -6817, 4235, 7191, -3600, -7511, 2934, 7769, -2247, -7969, 1541, 8104, -825, -8178, 101, 8186, 
--622, -8132, -1342, 8013, 2049, -7833, -2742, 7590, 3411, -7289, -4056, 6930, 4667, -6519, -5243, 6056, 5776, -5547, -6266, 4994, 6706, -4403, -7095, 3777, 7427, -3124, -7703, 2444, 7917, -1748, 
---8072, 1036, 8162, -319, -8191, -403, 8155, 1119, -8058, -1829, 7896, 2522, -7675, -3198, 7393, 3846, -7056, -4467, 6663, 5051, -6220, -5598, 5728, 6100, -5193, -6557, 4617, 6961, -4007, -7313, 
--3365, 7608, -2699, -7845, 2011, 8020, -1309, -8136, 595, 8187, 121, -8177, -838, 8103, 1546, -7969, -2244, 7772, 2923, -7517, -3581, 7203, 4210, -6836, -4809, 6414, 5368, -5946, -5889, 5431, 
--6362, -4877, -6789, 4283, 7161, -3659, -7482, 3005, 7743, -2331, -7947, 1637, 8089, -933, -8171, 220, 8189, 493, -8147, -1204, 8042, 1903, -7877, -2590, 7651, 3254, -7368, -3897, 7028, 4507, 
---6637, -5085, 6194, 5623, -5706, -6119, 5174, 6568, -4604, -6969, 3998, 7315, -3364, -7608, 2702, 7842, -2023, -8018, 1326, 8132, -622, -8187, -89, 8178, 797, -8110, -1501, 7979, 2191, -7791, 
---2867, 7541, 3519, -7238, -4146, 6878, 4741, -6469, -5301, 6009, 5820, -5507, -6297, 4961, 6725, -4381, -7104, 3766, 7429, -3126, -7700, 2460, 7911, -1778, -8066, 1080, 8158, -378, -8191, -330, 
--8162, 1033, -8074, -1730, 7924, 2412, -7717, -3078, 7451, 3719, -7131, -4334, 6757, 4915, -6335, -5461, 5864, 5965, -5352, -6426, 4799, 6838, -4212, -7201, 3592, 7508, -2947, -7763, 2279, 7957, 
---1597, -8096, 901, 8172, -200, -8190, -503, 8146, 1201, -8044, -1892, 7881, 2567, -7661, -3225, 7384, 3857, -7055, -4462, 6671, 5032, -6241, -5568, 5764, 6060, -5246, -6510, 4688, 6910, -4098, 
---7262, 3476, 7558, -2831, -7801, 2163, 7985, -1482, -8112, 788, 8179, -90, -8187, -609, 8134, 1303, -8024, -1988, 7854, 2657, -7628, -3309, 7345, 3934, -7010, -4532, 6623, 5096, -6190, -5624, 
--5710, 6109, -5191, -6552, 4632, 6946, -4042, -7290, 3421, 7580, -2777, -7818, 2112, 7996, -1433, -8119, 742, 8181, -48, -8186, -648, 8130, 1337, -8017, -2019, 7845, 2684, -7618, -3331, 7335, 
--3952, -7001, -4546, 6614, 5106, -6183, -5631, 5705, 6113, -5188, -6554, 4632, 6945, -4045, -7288, 3427, 7577, -2787, -7814, 2125, 7993, -1450, -8116, 763, 8180, -73, -8187, -620, 8134, 1306, 
---8024, -1984, 7856, 2646, -7634, -3291, 7355, 3911, -7026, -4504, 6645, 5064, -6219, -5589, 5747, 6072, -5237, -6514, 4687, 6908, -4106, -7255, 3495, 7548, -2860, -7790, 2204, 7974, -1534, -8104, 
--852, 8175, -166, -8190, -524, 8145, 1207, -8044, -1884, 7885, 2545, -7672, -3190, 7404, 3810, -7085, -4405, 6714, 4968, -6299, -5497, 5837, 5985, -5336, -6433, 4797, 6834, -4225, -7189, 3622, 
--7491, -2996, -7743, 2347, 7938, -1684, -8080, 1007, 8163, -325, -8191, -360, 8160, 1041, -8074, -1717, 7930, 2378, -7732, -3025, 7479, 3648, -7175, -4248, 6820, 4816, -6419, -5352, 5972, 5849, 
---5485, -6307, 4959, 6720, -4400, -7087, 3809, 7403, -3193, -7670, 2554, 7882, -1899, -8041, 1229, 8142, -552, -8189, -129, 8177, 808, -8111, -1483, 7987, 2146, -7809, -2795, 7576, 3423, -7293, 
---4030, 6958, 4606, -6577, -5153, 6148, 5661, -5680, -6133, 5170, 6561, -4628, -6945, 4051, 7280, -3449, -7567, 2822, 7799, -2177, -7980, 1516, 8105, -846, -8176, 169, 8189, 507, -8148, -1181, 
--8049, 1846, -7898, -2499, 7690, 3133, -7433, -3748, 7122, 4335, -6766, -4894, 6361, 5417, -5915, -5906, 5427, 6353, -4904, -6758, 4347, 7115, -3761, -7426, 3149, 7684, -2517, -7892, 1867, 8045, 
---1206, -8145, 535, 8188, 138, -8178, -811, 8110, 1477, -7990, -2134, 7813, 2775, -7587, -3399, 7307, 3998, -6979, -4571, 6603, 5112, -6185, -5620, 5723, 6089, -5225, -6518, 4690, 6901, -4125, 
---7240, 3531, 7528, -2916, -7768, 2279, 7954, -1629, -8088, 966, 8166, -299, -8191, -372, 8160, 1038, -8076, -1699, 7937, 2346, -7746, -2980, 7502, 3591, -7209, -4180, 6867, 4740, -6482, -5270, 
--6051, 5762, -5582, -6218, 5074, 6631, -4535, -7001, 3963, 7323, -3368, -7598, 2748, 7821, -2113, -7994, 1461, 8112, -802, -8178, 136, 8188, 528, -8146, -1191, 8048, 1844, -7900, -2487, 7697, 
--3111, -7445, -3716, 7142, 4295, -6795, -4847, 6401, 5365, -5967, -5850, 5491, 6294, -4982, -6699, 4439, 7057, -3868, -7372, 3270, 7635, -2653, -7851, 2017, 8013, -1369, -8125, 711, 8182, -51, 
---8187, -612, 8136, 1269, -8035, -1919, 7879, 2554, -7674, -3174, 7416, 3772, -7113, -4347, 6761, 4891, -6368, -5406, 5931, 5883, -5458, -6324, 4947, 6721, -4407, -7077, 3836, 7385, -3242, -7647, 
--2626, 7857, -1995, -8019, 1349, 8126, -696, -8183, 38, 8185, 619, -8137, -1274, 8033, 1918, -7880, -2552, 7674, 3167, -7421, -3763, 7118, 4333, -6772, -4877, 6380, 5388, -5949, -5865, 5478, 
--6303, -4974, -6703, 4436, 7057, -3872, -7368, 3282, 7629, -2672, -7844, 2044, 8007, -1404, -8120, 754, 8179, -102, -8188, -553, 8143, 1203, -8048, -1846, 7900, 2476, -7703, -3092, 7456, 3685, 
---7163, -4258, 6822, 4800, -6440, -5315, 6016, 5793, -5555, -6237, 5058, 6638, -4530, -7000, 3972, 7315, -3391, -7586, 2787, 7806, -2167, -7980, 1532, 8100, -889, -8172, 239, 8190, 411, -8158, 
---1060, 8073, 1699, -7939, -2330, 7754, 2945, -7521, -3542, 7239, 4115, -6914, -4664, 6543, 5181, -6134, -5668, 5684, 6117, -5201, -6530, 4683, 6899, -4138, -7228, 3565, 7509, -2973, -7745, 2359, 
--7930, -1734, -8068, 1095, 8154, -452, -8190, -195, 8174, 840, -8109, -1480, 7991, 2110, -7826, -2728, 7610, 3327, -7348, -3907, 7040, 4460, -6689, -4988, 6295, 5483, -5865, -5946, 5396, 6369, 
---4896, -6755, 4363, 7097, -3806, -7398, 3224, 7650, -2624, -7857, 2005, 8014, -1377, -8123, 738, 8180, -97, -8188, -546, 8145, 1184, -8053, -1816, 7909, 2435, -7719, -3041, 7480, 3626, -7197, 
---4191, 6868, 4728, -6499, -5237, 6088, 5713, -5642, -6155, 5160, 6558, -4648, -6922, 4106, 7242, -3541, -7519, 2953, 7749, -2349, -7933, 1728, 8067, -1100, -8154, 463, 8189, 175, -8177, -813, 
--8112, 1445, -8001, -2069, 7838, 2679, -7631, -3274, 7375, 3847, -7076, -4399, 6733, 4922, -6351, -5417, 5929, 5877, -5473, -6303, 4982, 6689, -4464, -7037, 3916, 7340, -3347, -7601, 2756, 7814, 
---2151, -7982, 1531, 8099, -904, -8170, 269, 8190, 364, -8163, -998, 8085, 1623, -7960, -2240, 7786, 2842, -7567, -3428, 7301, 3992, -6993, -4534, 6641, 5046, -6252, -5531, 5824, 5980, -5363, 
---6395, 4868, 6770, -4346, -7106, 3797, 7398, -3227, -7648, 2636, 7850, -2032, -8008, 1414, 8116, -790, -8178, 159, 8189, 471, -8154, -1100, 8068, 1720, -7937, -2331, 7756, 2927, -7532, -3507, 
--7262, 4064, -6950, -4599, 6596, 5105, -6205, -5582, 5776, 6025, -5314, -6433, 4819, 6802, -4299, -7133, 3751, 7419, -3183, -7664, 2595, 7862, -1993, -8016, 1378, 8120, -758, -8179, 131, 8188, 
--495, -8152, -1119, 8065, 1735, -7933, -2342, 7753, 2934, -7530, -3510, 7261, 4064, -6952, -4595, 6600, 5098, -6212, -5573, 5786, 6013, -5328, -6421, 4838, 6788, -4321, -7119, 3778, 7406, -3215, 
---7651, 2631, 7851, -2035, -8007, 1425, 8114, -808, -8176, 186, 8190, 436, -8157, -1057, 8076, 1670, -7950, -2274, 7777, 2864, -7560, -3439, 7298, 3991, -6996, -4523, 6652, 5026, -6272, -5503, 
--5854, 5946, -5405, -6356, 4922, 6728, -4414, -7063, 3878, 7355, -3323, -7608, 2746, 7815, -2156, -7979, 1552, 8095, -941, -8167, 323, 8190, 294, -8169, -912, 8099, 1523, -7985, -2126, 7824, 
--2715, -7620, -3291, 7371, 3846, -7082, -4380, 6751, 4888, -6384, -5370, 5979, 5819, -5542, -6237, 5071, 6617, -4575, -6963, 4050, 7266, -3505, -7531, 2938, 7750, -2357, -7928, 1760, 8060, -1156, 
---8147, 543, 8187, 70, -8183, -685, 8130, 1293, -8034, -1897, 7891, 2487, -7706, -3065, 7475, 3624, -7205, -4165, 6892, 4679, -6543, -5170, 6155, 5629, -5735, -6059, 5281, 6453, -4800, -6813, 
--4290, 7132, -3759, -7414, 3204, 7652, -2634, -7849, 2047, 8001, -1451, -8110, 846, 8173, -237, -8191, -374, 8162, 981, -8090, -1584, 7971, 2177, -7810, -2759, 7604, 3324, -7358, -3872, 7069, 
--4397, -6743, -4899, 6378, 5372, -5980, -5817, 5547, 6228, -5086, -6606, 4594, 6946, -4080, -7250, 3541, 7511, -2985, -7734, 2411, 7911, -1826, -8048, 1229, 8138, -627, -8185, 20, 8186, 585, 
---8143, -1188, 8055, 1783, -7924, -2369, 7748, 2941, -7531, -3498, 7272, 4034, -6975, -4550, 6638, 5039, -6267, -5503, 5860, 5934, -5424, -6335, 4956, 6699, -4463, -7029, 3944, 7319, -3406, -7570, 
--2848, 7779, -2276, -7948, 1690, 8071, -1097, -8153, 497, 8188, 104, -8181, -706, 8129, 1302, -8034, -1893, 7894, 2472, -7714, -3039, 7490, 3587, -7227, -4118, 6924, 4625, -6586, -5109, 6211, 
--5563, -5805, -5989, 5365, 6381, -4899, -6740, 4405, 7062, -3889, -7347, 3351, 7591, -2797, -7797, 2226, 7958, -1645, -8079, 1054, 8155, -460, -8190, -139, 8179, 735, -8126, -1328, 8028, 1913, 
---7890, -2489, 7707, 3050, -7486, -3596, 7223, 4121, -6924, -4626, 6587, 5104, -6216, -5558, 5811, 5979, -5377, -6371, 4913, 6727, -4425, -7050, 3912, 7333, -3381, -7579, 2829, 7784, -2265, -7949, 
--1688, 8071, -1103, -8152, 512, 8188, 81, -8183, -675, 8133, 1263, -8042, -1846, 7908, 2417, -7734, -2978, 7518, 3521, -7264, -4047, 6970, 4550, -6642, -5031, 6278, 5483, -5883, -5909, 5455, 
--6302, -5002, -6664, 4520, 6989, -4017, -7279, 3491, 7530, -2949, -7744, 2390, 7915, -1821, -8047, 1241, 8135, -656, -8184, 66, 8187, 522, -8151, -1109, 8070, 1688, -7950, -2260, 7786, 2819, 
---7585, -3364, 7342, 3890, -7064, -4398, 6748, 4881, -6398, -5341, 6014, 5771, -5602, -6174, 5158, 6542, -4691, -6879, 4197, 7179, -3684, -7444, 3151, 7668, -2603, -7855, 2040, 8000, -1469, -8106, 
--889, 8169, -306, -8191, -280, 8171, 862, -8110, -1442, 8006, 2012, -7864, -2574, 7679, 3120, -7458, -3653, 7196, 4164, -6901, -4657, 6568, 5124, -6204, -5566, 5807, 5978, -5383, -6362, 4930, 
--6712, -4453, -7029, 3953, 7309, -3435, -7554, 2897, 7759, -2347, -7926, 1784, 8052, -1213, -8139, 635, 8183, -56, -8188, -525, 8150, 1102, -8073, -1674, 7953, 2237, -7796, -2789, 7598, 3326, 
---7363, -3848, 7090, 4348, -6784, -4829, 6442, 5283, -6069, -5712, 5665, 6111, -5234, -6482, 4776, 6818, -4296, -7122, 3793, 7388, -3273, -7620, 2735, 7812, -2185, -7967, 1623, 8080, -1055, -8155, 
--480, 8188, 95, -8183, -671, 8134, 1242, -8048, -1809, 7920, 2364, -7755, -2910, 7550, 3439, -7309, -3953, 7031, 4445, -6720, -4918, 6374, 5364, -5999, -5785, 5593, 6176, -5161, -6538, 4702, 
--6867, -4222, -7163, 3720, 7423, -3202, -7647, 2666, 7833, -2119, -7982, 1560, 8090, -996, -8161, 425, 8189, 146, -8180, -718, 8129, 1284, -8040, -1845, 7911, 2396, -7745, -2937, 7539, 3461, 
---7299, -3970, 7022, 4458, -6712, -4926, 6368, 5369, -5996, -5787, 5593, 6174, -5164, -6534, 4709, 6861, -4234, -7156, 3736, 7414, -3222, -7639, 2691, 7824, -2149, -7974, 1595, 8084, -1036, -8157, 
--469, 8188, 97, -8183, -664, 8136, 1227, -8052, -1785, 7927, 2332, -7767, -2870, 7567, 3393, -7334, -3900, 7064, 4387, -6761, -4855, 6425, 5298, -6061, -5717, 5665, 6107, -5245, -6470, 4798, 
--6799, -4330, -7099, 3840, 7362, -3334, -7593, 2810, 7785, -2275, -7943, 1728, 8061, -1174, -8143, 613, 8184, -52, -8188, -512, 8152, 1071, -8080, -1626, 7967, 2172, -7819, -2710, 7632, 3232, 
---7411, -3741, 7154, 4231, -6865, -4702, 6542, 5149, -6190, -5574, 5808, 5971, -5400, -6341, 4965, 6680, -4509, -6989, 4031, 7264, -3535, -7506, 3021, 7711, -2496, -7883, 1957, 8015, -1411, -8113, 
--856, 8170, -300, -8191, -259, 8173, 815, -8118, -1369, 8024, 1915, -7895, -2453, 7727, 2978, -7525, -3491, 7287, 3985, -7017, -4463, 6712, 4918, -6379, -5353, 6015, 5760, -5625, -6143, 5207, 
--6495, -4767, -6820, 4304, 7110, -3822, -7371, 3322, 7595, -2808, -7786, 2280, 7939, -1744, -8058, 1197, 8138, -648, -8183, 93, 8188, 459, -8158, -1012, 8089, 1557, -7985, -2097, 7842, 2626, 
---7666, -3144, 7453, 3646, -7208, -4133, 6928, 4599, -6619, -5046, 6278, 5468, -5911, -5867, 5515, 6237, -5096, -6581, 4652, 6893, -4190, -7176, 3706, 7424, -3208, -7641, 2694, 7821, -2170, -7967, 
--1634, 8076, -1093, -8150, 545, 8186, 3, -8187, -553, 8149, 1098, -8076, -1640, 7965, 2172, -7821, -2697, 7639, 3207, -7426, -3705, 7177, 4184, -6898, -4646, 6587, 5085, -6248, -5503, 5880, 
--5895, -5487, -6262, 5068, 6599, -4629, -6909, 4167, 7186, -3689, -7433, 3193, 7645, -2684, -7824, 2162, 7967, -1633, -8077, 1094, 8149, -553, -8187, 8, 8186, 535, -8152, -1078, 8079, 1614, 
---7973, -2144, 7830, 2663, -7654, -3172, 7442, 3664, -7200, -4143, 6925, 4601, -6621, -5040, 6286, 5456, -5926, -5849, 5538, 6215, -5127, -6555, 4693, 6864, -4240, -7145, 3767, 7393, -3279, -7611, 
--2775, 7793, -2262, -7944, 1736, 8057, -1206, -8138, 668, 8181, -130, -8190, -411, 8162, 948, -8101, -1482, 8002, 2008, -7871, -2527, 7704, 3033, -7505, -3528, 7272, 4005, -7010, -4466, 6715, 
--4907, -6394, -5328, 6043, 5723, -5669, -6096, 5268, 6441, -4846, -6760, 4402, 7047, -3941, -7306, 3462, 7532, -2969, -7728, 2463, 7888, -1947, -8016, 1422, 8108, -893, -8168, 358, 8190, 176, 
---8179, -712, 8132, 1242, -8052, -1768, 7936, 2285, -7787, -2794, 7604, 3289, -7391, -3771, 7144, 4236, -6869, -4684, 6563, 5110, -6232, -5517, 5872, 5898, -5489, -6256, 5081, 6585, -4654, -6889, 
--4206, 7161, -3742, -7405, 3260, 7615, -2767, -7796, 2260, 7942, -1746, -8056, 1223, 8134, -697, -8180, 166, 8190, 364, -8167, -893, 8109, 1417, -8018, -1937, 7892, 2446, -7734, -2947, 7543, 
--3433, -7322, -3907, 7069, 4363, -6788, -4802, 6478, 5219, -6142, -5616, 5779, 5987, -5394, -6336, 4985, 6656, -4557, -6950, 4109, 7214, -3645, -7449, 3165, 7652, -2674, -7825, 2170, 7963, -1659, 
---8071, 1140, 8143, -618, -8184, 92, 8189, 433, -8162, -957, 8100, 1476, -8006, -1990, 7877, 2494, -7719, -2989, 7526, 3470, -7305, -3938, 7052, 4388, -6773, -4823, 6463, 5235, -6130, -5627, 
--5769, 5995, -5387, -6340, 4982, 6657, -4558, -6949, 4113, 7210, -3655, -7444, 3179, 7646, -2693, -7818, 2194, 7957, -1688, -8065, 1174, 8139, -657, -8182, 136, 8190, 384, -8166, -904, 8108, 
--1418, -8019, -1928, 7895, 2428, -7742, -2921, 7556, 3399, -7341, -3865, 7095, 4314, -6823, -4747, 6521, 5160, -6195, -5553, 5843, 5922, -5469, -6268, 5072, 6588, -4656, -6884, 4220, 7149, -3769, 
---7388, 3302, 7596, -2823, -7775, 2332, 7921, -1833, -8038, 1325, 8120, -814, -8173, 298, 8190, 217, -8178, -733, 8131, 1243, -8053, -1751, 7942, 2250, -7802, -2741, 7629, 3219, -7427, -3687, 
--7195, 4138, -6936, -4574, 6648, 4990, -6336, -5389, 5997, 5764, -5637, -6118, 5252, 6446, -4849, -6751, 4426, 7027, -3987, -7277, 3531, 7497, -3063, -7690, 2581, 7850, -2091, -7982, 1592, 8080, 
---1088, -8149, 579, 8184, -69, -8189, -443, 8161, 951, -8102, -1457, 8011, 1955, -7890, -2447, 7737, 2928, -7555, -3399, 7343, 3855, -7104, -4298, 6836, 4721, -6544, -5129, 6224, 5515, -5882, 
---5881, 5516, 6222, -5131, -6541, 4725, 6833, -4302, -7101, 3861, 7339, -3407, -7551, 2938, 7732, -2461, -7886, 1972, 8007, -1478, -8099, 976, 8158, -473, -8189, -34, 8185, 539, -8153, -1043, 
--8088, 1541, -7994, -2036, 7867, 2520, -7713, -2996, 7527, 3459, -7315, -3910, 7073, 4345, -6807, -4765, 6513, 5165, -6196, -5547, 5854, 5905, -5492, -6244, 5107, 6557, -4706, -6846, 4284, 7108, 
---3849, -7346, 3398, 7553, -2936, -7734, 2461, 7884, -1978, -8006, 1487, 8096, -993, -8158, 492, 8187, 7, -8187, -509, 8155, 1007, -8095, -1502, 8002, 1990, -7882, -2472, 7730, 2943, -7551, 
---3404, 7342, 3851, -7109, -4285, 6847, 4702, -6561, -5102, 6249, 5482, -5917, -5843, 5560, 6180, -5185, -6496, 4789, 6787, -4378, -7054, 3948, 7292, -3507, -7506, 3050, 7690, -2584, -7848, 2107, 
--7975, -1625, -8074, 1134, 8142, -642, -8182, 146, 8190, 349, -8170, -845, 8118, 1335, -8038, -1822, 7927, 2300, -7789, -2771, 7620, 3230, -7426, -3680, 7203, 4113, -6956, -4534, 6682, 4936, 
---6385, -5322, 6064, 5686, -5722, -6032, 5358, 6353, -4977, -6654, 4575, 6928, -4160, -7179, 3727, 7402, -3283, -7600, 2826, 7769, -2360, -7911, 1885, 8024, -1404, -8109, 917, 8163, -429, -8189, 
---63, 8185, 552, -8153, -1041, 8089, 1525, -7999, -2004, 7878, 2474, -7731, -2937, 7555, 3388, -7353, -3828, 7124, 4252, -6871, -4663, 6592, 5056, -6291, -5432, 5966, 5786, -5622, -6122, 5257, 
--6435, -4875, -6726, 4473, 6991, -4058, -7233, 3627, 7448, -3185, -7638, 2730, 7800, -2268, -7935, 1796, 8041, -1319, -8120, 837, 8169, -353, -8191, -133, 8182, 617, -8146, -1101, 8080, 1578, 
---7988, -2052, 7865, 2516, -7717, -2974, 7541, 3418, -7340, -3853, 7111, 4272, -6860, -4678, 6582, 5066, -6285, -5437, 5963, 5788, -5623, -6121, 5261, 6430, -4883, -6718, 4487, 6981, -4077, -7222, 
--3651, 7436, -3214, -7626, 2765, 7787, -2308, -7924, 1842, 8031, -1371, -8113, 894, 8164, -416, -8190, -65, 8185, 544, -8154, -1023, 8093, 1496, -8006, -1966, 7890, 2426, -7749, -2881, 7580, 
--3323, -7387, -3756, 7166, 4174, -6923, -4579, 6655, 4966, -6366, -5339, 6054, 5691, -5723, -6026, 5370, 6338, -5002, -6630, 4615, 6898, -4214, -7144, 3797, 7364, -3370, -7561, 2929, 7731, -2481, 
---7876, 2022, 7992, -1559, -8084, 1089, 8146, -617, -8183, 141, 8190, 333, -8172, -807, 8124, 1277, -8051, -1744, 7949, 2203, -7822, -2657, 7668, 3099, -7489, -3533, 7284, 3953, -7057, -4362, 
--6804, 4754, -6530, -5132, 6233, 5491, -5918, -5833, 5580, 6154, -5227, -6456, 4854, 6734, -4467, -6992, 4063, 7225, -3649, -7436, 3220, 7620, -2783, -7781, 2335, 7914, -1881, -8023, 1419, 8104, 
---955, -8160, 486, 8187, -18, -8189, -453, 8162, 920, -8110, -1385, 8030, 1844, -7925, -2298, 7793, 2743, -7637, -3181, 7454, 3606, -7249, -4021, 7018, 4421, -6767, -4808, 6491, 5177, -6197, 
---5532, 5881, 5866, -5547, -6183, 5194, 6478, -4826, -6754, 4441, 7006, -4043, -7237, 3630, 7442, -3208, -7625, 2774, 7782, -2333, -7915, 1882, 8021, -1428, -8103, 967, 8157, -506, -8187, 41, 
--8188, 422, -8165, -886, 8114, 1344, -8039, -1800, 7936, 2248, -7810, -2691, 7657, 3122, -7482, -3546, 7280, 3956, -7058, -4355, 6811, 4739, -6545, -5109, 6256, 5461, -5949, -5797, 5621, 6112, 
---5278, -6411, 4916, 6686, -4541, -6943, 4150, 7175, -3747, -7387, 3331, 7573, -2907, -7737, 2472, 7875, -2031, -7990, 1581, 8077, -1129, -8142, 672, 8178, -215, -8191, -245, 8177, 702, -8139, 
---1158, 8073, 1608, -7984, -2056, 7868, 2494, -7730, -2927, 7565, 3349, -7379, -3761, 7168, 4160, -6937, -4548, 6683, 4920, -6410, -5278, 6115, 5617, -5803, -5941, 5471, 6245, -5125, -6531, 4761, 
--6794, -4384, -7039, 3992, 7260, -3590, -7460, 3175, 7635, -2752, -7789, 2319, 7916, -1881, -8022, 1436, 8100, -988, -8156, 536, 8185, -84, -8190, -370, 8169, 821, -8124, -1271, 8053, 1715, 
---7959, -2155, 7840, 2587, -7698, -3013, 7531, 3427, -7343, -3833, 7130, 4225, -6899, -4605, 6644, 4970, -6372, -5322, 6078, 5655, -5768, -5973, 5439, 6271, -5095, -6552, 4734, 6811, -4361, -7051, 
--3973, 7268, -3576, -7465, 3165, 7638, -2748, -7789, 2320, 7915, -1888, -8020, 1448, 8098, -1006, -8154, 559, 8184, -113, -8191, -336, 8171, 781, -8130, -1225, 8062, 1664, -7972, -2100, 7857, 
--2527, -7720, -2949, 7558, 3360, -7376, -3762, 7171, 4151, -6946, -4530, 6698, 4893, -6433, -5244, 6148, 5577, -5846, -5895, 5525, 6194, -5190, -6476, 4837, 6738, -4473, -6981, 4094, 7202, -3705, 
---7404, 3303, 7581, -2894, -7739, 2474, 7872, -2050, -7984, 1617, 8070, -1182, -8135, 742, 8174, -302, -8191, -141, 8183, 581, -8152, -1021, 8096, 1457, -8019, -1889, 7916, 2315, -7792, -2735, 
--7644, 3145, -7476, -3548, 7285, 3938, -7074, -4319, 6841, 4685, -6591, -5040, 6319, 5378, -6032, -5702, 5725, 6008, -5405, -6298, 5066, 6569, -4716, -6822, 4350, 7054, -3974, -7267, 3584, 7458, 
---3187, -7629, 2778, 7776, -2364, -7903, 1942, 8006, -1516, -8088, 1083, 8144, -650, -8180, 214, 8190, 221, -8180, -657, 8144, 1090, -8087, -1520, 8005, 1945, -7903, -2366, 7776, 2777, -7630, 
---3183, 7460, 3578, -7271, -3964, 7060, 4338, -6831, -4700, 6581, 5048, -6315, -5383, 6029, 5701, -5729, -6005, 5410, 6290, -5079, -6559, 4731, 6808, -4373, -7040, 4001, 7250, -3619, -7442, 3226, 
--7611, -2826, -7761, 2416, 7887, -2002, -7993, 1580, 8075, -1157, -8137, 728, 8174, -299, -8191, -132, 8183, 561, -8155, -990, 8102, 1414, -8029, -1835, 7931, 2250, -7815, -2660, 7674, 3061, 
---7515, -3456, 7333, 3838, -7134, -4212, 6912, 4572, -6674, -4922, 6416, 5256, -6143, -5578, 5851, 5882, -5545, -6172, 5223, 6443, -4888, -6699, 4538, 6934, -4178, -7152, 3805, 7349, -3424, -7528, 
--3031, 7685, -2633, -7823, 2226, 7937, -1815, -8032, 1397, 8104, -978, -8156, 554, 8183, -131, -8191, -294, 8175, 717, -8139, -1139, 8079, 1556, -7999, -1970, 7897, 2377, -7775, -2780, 7630, 
--3173, -7468, -3559, 7283, 3934, -7081, -4300, 6859, 4652, -6620, -4994, 6362, 5320, -6089, -5635, 5798, 5932, -5494, -6215, 5174, 6480, -4842, -6730, 4495, 6960, -4139, -7173, 3770, 7365, -3393, 
---7540, 3006, 7693, -2613, -7828, 2211, 7940, -1806, -8034, 1394, 8104, -980, -8155, 563, 8183, -146, -8191, -274, 8176, 690, -8142, -1106, 8085, 1518, -8008, -1927, 7909, 2329, -7792, -2726, 
--7652, 3115, -7494, -3497, 7316, 3868, -7120, -4231, 6904, 4580, -6672, -4920, 6422, 5245, -6157, -5558, 5874, 5855, -5578, -6139, 5266, 6404, -4943, -6655, 4605, 6888, -4257, -7104, 3897, 7300, 
---3529, -7479, 3150, 7637, -2766, -7778, 2372, 7897, -1975, -7997, 1571, 8075, -1165, -8135, 754, 8172, -344, -8190, -70, 8186, 480, -8163, -892, 8117, 1299, -8053, -1704, 7966, 2103, -7862, 
---2499, 7735, 2886, -7591, -3267, 7427, 3638, -7245, -4002, 7044, 4354, -6827, -4696, 6591, 5025, -6341, -5343, 6073, 5645, -5792, -5936, 5495, 6209, -5186, -6469, 4862, 6710, -4529, -6937, 4182, 
--7144, -3827, -7336, 3461, 7507, -3088, -7662, 2706, 7795, -2320, -7911, 1926, 8006, -1529, -8083, 1127, 8138, -724, -8175, 318, 8190, 87, -8186, -494, 8161, 897, -8117, -1300, 8052, 1697, 
---7969, -2092, 7865, 2480, -7743, -2863, 7601, 3238, -7442, -3606, 7263, 3963, -7069, -4313, 6855, 4649, -6627, -4977, 6381, 5290, -6122, -5592, 5846, 5879, -5558, -6153, 5254, 6410, -4940, -6654, 
--4613, 6879, -4276, -7090, 3927, 7281, -3571, -7457, 3205, 7613, -2833, -7753, 2453, 7872, -2068, -7974, 1677, 8055, -1285, -8119, 887, 8162, -489, -8186, 89, 8190, 310, -8176, -709, 8140, 
--1105, -8087, -1500, 8013, 1889, -7922, -2276, 7810, 2655, -7682, -3029, 7534, 3394, -7370, -3753, 7187, 4101, -6989, -4441, 6773, 4769, -6542, -5087, 6295, 5391, -6035, -5684, 5759, 5962, -5471, 
---6227, 5169, 6476, -4857, -6712, 4532, 6930, -4198, -7134, 3853, 7319, -3500, -7488, 3138, 7639, -2771, -7773, 2396, 7888, -2017, -7986, 1632, 8063, -1245, -8124, 853, 8164, -462, -8187, 68, 
--8189, 324, -8175, -717, 8140, 1107, -8087, -1495, 8015, 1878, -7926, -2259, 7817, 2632, -7692, -3001, 7547, 3361, -7388, -3715, 7209, 4058, -7016, -4394, 6806, 4718, -6582, -5033, 6341, 5334, 
---6087, -5625, 5819, 5901, -5539, -6166, 5244, 6414, -4940, -6650, 4623, 6869, -4298, -7074, 3961, 7261, -3617, -7433, 3264, 7587, -2905, -7726, 2538, 7845, -2167, -7949, 1790, 8033, -1411, -8100, 
--1027, 8148, -643, -8179, 255, 8190, 131, -8185, -518, 8160, 902, -8118, -1286, 8057, 1664, -7979, -2041, 7882, 2411, -7770, -2778, 7638, 3136, -7491, -3489, 7326, 3832, -7147, -4169, 6951, 
--4494, -6741, -4811, 6514, 5116, -6275, -5411, 6021, 5692, -5755, -5962, 5475, 6217, -5186, -6461, 4883, 6688, -4571, -6903, 4248, 7100, -3917, -7284, 3576, 7450, -3230, -7601, 2875, 7734, -2515, 
---7852, 2149, 7951, -1780, -8035, 1405, 8099, -1030, -8148, 650, 8178, -271, -8191, -110, 8185, 489, -8163, -868, 8122, 1244, -8065, -1618, 7990, 1987, -7899, -2354, 7789, 2713, -7664, -3068, 
--7522, 3415, -7365, -3756, 7190, 4086, -7003, -4410, 6798, 4723, -6582, -5027, 6349, 5319, -6105, -5601, 5847, 5869, -5578, -6126, 5295, 6368, -5003, -6599, 4699, 6814, -4388, -7016, 4065, 7202, 
---3736, -7374, 3397, 7529, -3053, -7669, 2701, 7792, -2345, -7900, 1983, 7990, -1619, -8065, 1249, 8121, -880, -8162, 506, 8184, -134, -8191, -241, 8179, 612, -8152, -985, 8107, 1352, -8046, 
---1719, 7967, 2081, -7873, -2439, 7762, 2791, -7636, -3139, 7492, 3478, -7336, -3811, 7162, 4135, -6976, -4452, 6773, 4757, -6559, -5055, 6329, 5340, -6088, -5617, 5834, 5879, -5569, -6132, 5291, 
--6369, -5005, -6596, 4707, 6807, -4401, -7007, 4084, 7190, -3761, -7360, 3429, 7513, -3092, -7653, 2747, 7776, -2399, -7884, 2044, 7975, -1687, -8052, 1325, 8110, -963, -8154, 596, 8180, -231, 
---8191, -137, 8184, 502, -8163, -868, 8123, 1230, -8069, -1591, 7997, 1947, -7911, -2301, 7808, 2648, -7691, -2992, 7556, 3327, -7409, -3658, 7245, 3979, -7069, -4295, 6877, 4599, -6674, -4897, 
--6456, 5183, -6227, -5460, 5983, 5724, -5731, -5979, 5465, 6220, -5190, -6451, 4904, 6667, -4610, -6872, 4305, 7061, -3994, -7239, 3673, 7400, -3347, -7549, 3013, 7680, -2676, -7799, 2331, 7901, 
---1984, -7989, 1631, 8060, -1278, -8117, 920, 8157, -562, -8183, 202, 8190, 157, -8185, -517, 8161, 874, -8124, -1231, 8069, 1583, -8000, -1935, 7915, 2280, -7816, -2623, 7700, 2958, -7572, 
---3290, 7427, 3613, -7271, -3932, 7098, 4240, -6914, -4543, 6715, 4834, -6506, -5118, 6282, 5391, -6048, -5655, 5802, 5906, -5546, -6148, 5278, 6376, -5002, -6594, 4715, 6798, -4421, -6990, 4117, 
--7168, -3808, -7334, 3489, 7484, -3167, -7622, 2836, 7743, -2502, -7852, 2162, 7945, -1820, -8024, 1473, 8087, -1125, -8136, 774, 8169, -423, -8188, 70, 8190, 282, -8179, -635, 8150, 984, 
---8109, -1333, 8051, 1678, -7980, -2021, 7892, 2358, -7792, -2693, 7676, 3021, -7547, -3345, 7403, 3661, -7248, -3972, 7077, 4273, -6895, -4569, 6699, 4854, -6493, -5132, 6273, 5398, -6044, -5657, 
--5802, 5903, -5552, -6140, 5289, 6364, -5020, -6579, 4739, 6779, -4452, -6969, 4155, 7145, -3853, -7309, 3542, 7458, -3227, -7596, 2904, 7718, -2578, -7828, 2246, 7922, -1912, -8004, 1573, 8069, 
---1233, -8122, 889, 8159, -546, -8183, 200, 8190, 144, -8185, -490, 8164, 833, -8130, -1176, 8079, 1515, -8017, -1853, 7938, 2185, -7847, -2515, 7740, 2839, -7622, -3160, 7489, 3473, -7344, 
---3781, 7185, 4081, -7015, -4375, 6831, 4660, -6638, -4938, 6430, 5206, -6214, -5466, 5985, 5715, -5748, -5955, 5498, 6184, -5242, -6403, 4974, 6609, -4700, -6805, 4416, 6988, -4127, -7160, 3829, 
--7318, -3526, -7466, 3215, 7598, -2901, -7719, 2580, 7825, -2257, -7920, 1928, 7998, -1599, -8065, 1264, 8117, -930, -8156, 592, 8180, -255, -8191, -83, 8187, 420, -8170, -757, 8138, 1091, 
---8094, -1426, 8035, 1755, -7963, -2083, 7877, 2406, -7779, -2726, 7666, 3040, -7542, -3350, 7404, 3652, -7256, -3950, 7093, 4240, -6920, -4524, 6734, 4798, -6539, -5066, 6331, 5324, -6115, -5574, 
--5887, 5814, -5650, -6045, 5403, 6264, -5149, -6475, 4885, 6672, -4614, -6861, 4334, 7036, -4049, -7202, 3756, 7353, -3458, -7494, 3153, 7621, -2846, -7738, 2531, 7839, -2215, -7930, 1893, 8005, 
---1570, -8070, 1243, 8119, -916, -8157, 586, 8180, -257, -8191, -74, 8187, 403, -8172, -733, 8141, 1060, -8100, -1387, 8043, 1709, -7975, -2030, 7893, 2346, -7799, -2660, 7692, 2968, -7574, 
---3272, 7442, 3569, -7300, -3862, 7144, 4147, -6979, -4427, 6801, 4698, -6615, -4963, 6416, 5218, -6208, -5467, 5989, 5705, -5763, -5935, 5526, 6154, -5282, -6365, 5028, 6564, -4768, -6755, 4498, 
--6932, -4224, -7101, 3941, 7256, -3655, -7402, 3360, 7534, -3063, -7657, 2759, 7765, -2452, -7863, 2141, 7946, -1828, -8020, 1510, 8078, -1192, -8126, 871, 8160, -550, -8182, 227, 8190, 95, 
---8187, -418, 8170, 738, -8142, -1059, 8099, 1376, -8046, -1693, 7979, 2005, -7901, -2316, 7810, 2620, -7708, -2923, 7593, 3219, -7468, -3512, 7329, 3798, -7182, -4079, 7022, 4352, -6853, -4621, 
--6672, 4880, -6483, -5133, 6282, 5377, -6073, -5614, 5854, 5841, -5628, -6061, 5392, 6269, -5149, -6470, 4897, 6659, -4640, -6840, 4374, 7008, -4103, -7168, 3825, 7315, -3543, -7453, 3254, 7578, 
---2962, -7693, 2664, 7795, -2364, -7887, 2059, 7966, -1753, -8034, 1443, 8089, -1133, -8133, 819, 8164, -506, -8184, 190, 8190, 123, -8187, -438, 8169, 750, -8141, -1063, 8099, 1373, -8048, 
---1682, 7983, 1986, -7908, -2289, 7819, 2587, -7721, -2883, 7610, 3172, -7490, -3459, 7358, 3738, -7216, -4014, 7062, 4281, -6900, -4545, 6727, 4800, -6545, -5049, 6353, 5289, -6153, -5524, 5942, 
--5748, -5726, -5966, 5499, 6173, -5266, -6373, 5024, 6562, -4777, -6744, 4521, 6914, -4261, -7075, 3993, 7225, -3722, -7366, 3443, 7495, -3162, -7615, 2874, 7722, -2585, -7820, 2290, 7905, -1994, 
---7981, 1693, 8044, -1392, -8097, 1088, 8137, -784, -8167, 477, 8184, -172, -8191, -135, 8185, 440, -8170, -746, 8141, 1049, -8103, -1352, 8052, 1652, -7991, -1950, 7917, 2244, -7835, -2536, 
--7740, 2823, -7636, -3108, 7519, 3386, -7394, -3661, 7258, 3930, -7113, -4194, 6957, 4451, -6793, -4703, 6618, 4947, -6436, -5186, 6243, 5416, -6044, -5640, 5835, 5854, -5620, -6062, 5396, 6260, 
---5166, -6451, 4928, 6631, -4685, -6805, 4434, 6967, -4179, -7121, 3917, 7264, -3651, -7399, 3379, 7522, -3104, -7636, 2824, 7739, -2542, -7833, 2254, 7914, -1966, -7987, 1673, 8047, -1381, -8098, 
--1084, 8137, -789, -8166, 490, 8183, -194, -8191, -105, 8187, 402, -8173, -700, 8147, 994, -8111, -1290, 8064, 1581, -8007, -1872, 7939, 2159, -7861, -2444, 7772, 2724, -7675, -3002, 7565, 
--3274, -7448, -3544, 7319, 3807, -7183, -4067, 7035, 4319, -6881, -4568, 6716, 4808, -6544, -5045, 6362, 5272, -6173, -5495, 5975, 5708, -5771, -5916, 5558, 6114, -5341, -6306, 5114, 6488, -4883, 
---6664, 4644, 6828, -4401, -6987, 4151, 7134, -3897, -7274, 3637, 7402, -3374, -7523, 3106, 7633, -2835, -7735, 2559, 7825, -2282, -7907, 2001, 7977, -1719, -8038, 1433, 8088, -1147, -8130, 859, 
--8159, -571, -8180, 281, 8189, 8, -8190, -298, 8179, 585, -8159, -874, 8127, 1159, -8087, -1445, 8035, 1727, -7976, -2008, 7904, 2285, -7825, -2560, 7734, 2831, -7636, -3099, 7526, 3362, 
---7409, -3623, 7282, 3876, -7147, -4127, 7002, 4371, -6850, -4611, 6688, 4843, -6520, -5072, 6342, 5292, -6159, -5507, 5966, 5714, -5769, -5915, 5562, 6108, -5351, -6295, 5131, 6472, -4908, -6643, 
--4677, 6804, -4442, -6959, 4200, 7103, -3955, -7241, 3704, 7368, -3451, -7488, 3191, 7597, -2930, -7699, 2664, 7790, -2396, -7873, 2124, 7946, -1852, -8010, 1576, 8063, -1300, -8109, 1020, 8143, 
---742, -8169, 461, 8184, -181, -8191, -100, 8187, 379, -8175, -659, 8152, 937, -8120, -1215, 8078, 1490, -8028, -1764, 7967, 2035, -7899, -2305, 7819, 2570, -7733, -2833, 7636, 3092, -7532, 
---3348, 7417, 3599, -7296, -3847, 7165, 4089, -7027, -4328, 6880, 4559, -6727, -4788, 6564, 5009, -6396, -5225, 6219, 5434, -6036, -5639, 5846, 5834, -5650, -6026, 5446, 6208, -5239, -6385, 5023, 
--6552, -4804, -6715, 4578, 6867, -4349, -7014, 4113, 7151, -3874, -7281, 3630, 7402, -3384, -7516, 3132, 7619, -2878, -7716, 2620, 7803, -2361, -7882, 2097, 7951, -1834, -8013, 1566, 8064, -1299, 
---8108, 1029, 8142, -760, -8168, 488, 8183, -218, -8191, -54, 8188, 324, -8179, -596, 8158, 864, -8130, -1134, 8092, 1400, -8047, -1666, 7991, 1928, -7928, -2190, 7855, 2448, -7776, -2704, 
--7686, 2956, -7590, -3206, 7484, 3450, -7372, -3693, 7250, 3929, -7122, -4164, 6985, 4391, -6842, -4616, 6690, 4833, -6534, -5047, 6368, 5254, -6198, -5457, 6019, 5652, -5836, -5843, 5645, 6025, 
---5450, -6203, 5248, 6373, -5042, -6537, 4829, 6693, -4613, -6843, 4391, 6984, -4166, -7120, 3934, 7246, -3701, -7367, 3462, 7477, -3222, -7582, 2977, 7677, -2731, -7766, 2480, 7845, -2228, -7918, 
--1973, 7980, -1718, -8036, 1459, 8082, -1201, -8121, 939, 8150, -679, -8173, 417, 8185, -156, -8191, -106, 8187, 367, -8176, -629, 8155, 888, -8128, -1147, 8091, 1404, -8047, -1661, 7993, 
--1914, -7933, -2167, 7863, 2415, -7788, -2663, 7702, 2906, -7611, -3148, 7511, 3385, -7405, -3620, 7289, 3849, -7169, -4076, 7039, 4297, -6905, -4516, 6762, 4728, -6614, -4937, 6458, 5139, -6297, 
---5338, 6128, 5529, -5956, -5717, 5776, 5897, -5592, -6073, 5401, 6241, -5206, -6405, 5005, 6560, -4801, -6711, 4591, 6853, -4378, -6991, 4159, 7120, -3939, -7243, 3712, 7358, -3484, -7467, 3251, 
--7567, -3018, -7662, 2779, 7747, -2540, -7826, 2296, 7896, -2053, -7961, 1806, 8016, -1559, -8065, 1309, 8104, -1060, -8138, 808, 8162, -558, -8180, 305, 8189, -54, -8191, -198, 8184, 449, 
---8171, -701, 8149, 949, -8121, -1199, 8083, 1446, -8040, -1692, 7987, 1936, -7929, -2179, 7861, 2418, -7789, -2656, 7707, 2890, -7620, -3123, 7524, 3351, -7423, -3577, 7313, 3798, -7199, -4018, 
--7076, 4231, -6949, -4443, 6813, 4648, -6673, -4851, 6526, 5047, -6374, -5241, 6215, 5427, -6052, -5611, 5882, 5787, -5709, -5960, 5529, 6125, -5345, -6287, 5156, 6441, -4963, -6591, 4764, 6733, 
---4564, -6870, 4357, 7000, -4148, -7125, 3934, 7241, -3719, -7353, 3499, 7457, -3277, -7556, 3051, 7645, -2824, -7731, 2593, 7807, -2362, -7878, 2127, 7940, -1892, -7997, 1654, 8045, -1417, -8088, 
--1176, 8122, -937, -8151, 695, 8170, -455, -8185, 212, 8190, 29, -8190, -271, 8181, 511, -8167, -752, 8144, 990, -8116, -1230, 8079, 1466, -8037, -1703, 7986, 1936, -7930, -2169, 7866, 
--2398, -7797, -2627, 7719, 2851, -7637, -3075, 7546, 3294, -7451, -3512, 7348, 3725, -7240, -3936, 7125, 4142, -7006, -4347, 6878, 4545, -6748, -4742, 6609, 4932, -6467, -5121, 6318, 5302, -6166, 
---5481, 6007, 5654, -5845, -5823, 5676, 5986, -5504, -6145, 5327, 6298, -5146, -6447, 4960, 6588, -4772, -6726, 4578, 6856, -4383, -6983, 4182, 7102, -3979, -7216, 3772, 7323, -3564, -7426, 3351, 
--7521, -3137, -7611, 2920, 7693, -2702, -7771, 2480, 7840, -2258, -7906, 2032, 7962, -1807, -8015, 1579, 8058, -1352, -8098, 1122, 8128, -893, -8155, 661, 8172, -432, -8185, 200, 8190, 30, 
---8190, -261, 8182, 491, -8169, -721, 8148, 949, -8122, -1178, 8088, 1404, -8050, -1630, 8003, 1853, -7952, -2077, 7893, 2296, -7830, -2516, 7759, 2731, -7684, -2946, 7601, 3157, -7514, -3367, 
--7419, 3572, -7321, -3776, 7215, 3976, -7106, -4174, 6989, 4366, -6869, -4557, 6742, 4743, -6612, -4927, 6475, 5104, -6335, -5280, 6189, 5450, -6040, -5617, 5884, 5778, -5726, -5936, 5562, 6088, 
---5396, -6237, 5224, 6379, -5050, -6518, 4871, 6651, -4690, -6780, 4504, 6902, -4316, -7021, 4124, 7132, -3930, -7240, 3732, 7341, -3533, -7438, 3330, 7527, -3127, -7613, 2919, 7691, -2712, -7766, 
--2500, 7832, -2289, -7895, 2075, 7950, -1861, -8002, 1644, 8045, -1428, -8085, 1210, 8116, -992, -8144, 772, 8164, -554, -8179, 333, 8187, -115, -8191, -106, 8188, 324, -8180, -544, 8164, 
--761, -8145, -980, 8118, 1195, -8087, -1412, 8048, 1625, -8006, -1839, 7956, 2050, -7903, -2260, 7842, 2468, -7777, -2675, 7706, 2878, -7630, -3081, 7548, 3279, -7462, -3477, 7369, 3671, -7274, 
---3864, 7171, 4051, -7065, -4238, 6953, 4420, -6838, -4601, 6716, 4776, -6591, -4950, 6461, 5118, -6328, -5285, 6188, 5445, -6047, -5604, 5900, 5757, -5751, -5908, 5596, 6053, -5439, -6196, 5277, 
--6332, -5113, -6466, 4944, 6593, -4774, -6718, 4599, 6836, -4423, -6952, 4242, 7060, -4061, -7166, 3875, 7265, -3688, -7361, 3498, 7450, -3307, -7536, 3112, 7616, -2917, -7691, 2719, 7760, -2521, 
---7826, 2319, 7884, -2118, -7939, 1914, 7987, -1711, -8032, 1505, 8070, -1300, -8104, 1092, 8131, -886, -8154, 678, 8170, -471, -8183, 263, 8189, -56, -8191, -153, 8186, 359, -8178, -567, 
--8163, 772, -8145, -979, 8119, 1183, -8090, -1387, 8054, 1589, -8015, -1792, 7969, 1991, -7920, -2191, 7864, 2387, -7805, -2584, 7740, 2776, -7671, -2969, 7596, 3158, -7518, -3346, 7434, 3531, 
---7347, -3715, 7253, 3894, -7157, -4073, 7055, 4247, -6951, -4421, 6840, 4589, -6727, -4757, 6609, 4920, -6488, -5081, 6361, 5237, -6233, -5392, 6099, 5541, -5964, -5689, 5823, 5831, -5680, -5972, 
--5533, 6106, -5384, -6239, 5230, 6367, -5075, -6492, 4915, 6611, -4755, -6728, 4589, 6839, -4424, -6948, 4253, 7051, -4083, -7151, 3908, 7245, -3733, -7337, 3554, 7422, -3375, -7505, 3192, 7581, 
---3010, -7655, 2823, 7722, -2638, -7787, 2449, 7845, -2261, -7900, 2070, 7949, -1880, -7995, 1687, 8035, -1495, -8071, 1300, 8102, -1107, -8129, 911, 8150, -718, -8168, 521, 8180, -327, -8188, 
--131, 8190, 63, -8190, -259, 8183, 452, -8173, -647, 8157, 840, -8138, -1034, 8112, 1225, -8084, -1417, 8050, 1606, -8013, -1796, 7970, 1983, -7924, -2170, 7872, 2355, -7817, -2539, 7757, 
--2720, -7694, -2902, 7625, 3080, -7554, -3257, 7477, 3431, -7397, -3605, 7312, 3775, -7225, -3944, 7132, 4109, -7038, -4274, 6937, 4434, -6835, -4594, 6728, 4749, -6619, -4903, 6504, 5052, -6388, 
---5201, 6267, 5345, -6145, -5488, 6017, 5625, -5889, -5762, 5755, 5893, -5621, -6023, 5481, 6148, -5341, -6272, 5197, 6390, -5052, -6506, 4902, 6617, -4752, -6727, 4597, 6830, -4442, -6933, 4284, 
--7029, -4125, -7124, 3962, 7213, -3799, -7300, 3633, 7381, -3467, -7461, 3297, 7534, -3128, -7606, 2955, 7672, -2783, -7735, 2608, 7793, -2433, -7849, 2256, 7898, -2079, -7946, 1900, 7988, -1722, 
---8027, 1542, 8061, -1362, -8092, 1181, 8118, -1001, -8141, 818, 8158, -637, -8173, 455, 8182, -274, -8189, 91, 8190, 89, -8190, -272, 8183, 452, -8174, -633, 8159, 812, -8142, -993, 
--8119, 1171, -8094, -1350, 8063, 1526, -8031, -1703, 7992, 1877, -7952, -2052, 7906, 2224, -7859, -2397, 7805, 2567, -7750, -2736, 7690, 2903, -7628, -3070, 7560, 3233, -7491, -3397, 7416, 3557, 
---7340, -3717, 7258, 3873, -7176, -4029, 7088, 4181, -6998, -4333, 6904, 4480, -6809, -4628, 6708, 4771, -6607, -4914, 6500, 5052, -6393, -5190, 6281, 5324, -6168, -5456, 6050, 5585, -5932, -5712, 
--5809, 5835, -5686, -5957, 5559, 6074, -5431, -6190, 5298, 6302, -5166, -6412, 5029, 6517, -4892, -6622, 4751, 6721, -4611, -6819, 4466, 6912, -4321, -7004, 4173, 7091, -4025, -7176, 3874, 7257, 
---3723, -7335, 3568, 7409, -3414, -7481, 3257, 7548, -3101, -7614, 2941, 7674, -2782, -7733, 2621, 7787, -2460, -7839, 2297, 7885, -2134, -7930, 1969, 7970, -1806, -8008, 1639, 8041, -1474, -8073, 
--1307, 8098, -1142, -8123, 974, 8142, -808, -8159, 640, 8172, -473, -8182, 305, 8187, -139, -8191, -29, 8190, 195, -8187, -363, 8178, 528, -8169, -695, 8154, 859, -8137, -1025, 8115, 
--1188, -8092, -1353, 8064, 1514, -8035, -1677, 8000, 1837, -7964, -1998, 7923, 2157, -7880, -2316, 7833, 2472, -7784, -2628, 7731, 2782, -7676, -2936, 7617, 3087, -7556, -3238, 7491, 3387, -7424, 
---3535, 7353, 3680, -7281, -3825, 7204, 3967, -7127, -4109, 7045, 4247, -6962, -4385, 6875, 4520, -6787, -4654, 6694, 4785, -6601, -4915, 6504, 5042, -6406, -5168, 6304, 5290, -6201, -5413, 6095, 
--5530, -5988, -5648, 5877, 5762, -5766, -5875, 5651, 5983, -5536, -6092, 5417, 6195, -5298, -6299, 5175, 6398, -5053, -6496, 4926, 6590, -4800, -6684, 4671, 6772, -4542, -6861, 4409, 6944, -4277, 
---7027, 4142, 7105, -4007, -7183, 3869, 7256, -3732, -7328, 3591, 7395, -3451, -7461, 3309, 7523, -3167, -7584, 3022, 7641, -2879, -7696, 2732, 7747, -2587, -7796, 2439, 7841, -2293, -7885, 2144, 
--7925, -1996, -7963, 1846, 7997, -1697, -8029, 1546, 8057, -1396, -8084, 1244, 8107, -1094, -8128, 942, 8144, -792, -8160, 639, 8171, -489, -8181, 336, 8186, -186, -8191, 34, 8190, 116, 
---8189, -268, 8183, 417, -8177, -568, 8165, 717, -8153, -868, 8136, 1015, -8119, -1165, 8096, 1311, -8073, -1460, 8046, 1605, -8018, -1752, 7985, 1896, -7952, -2041, 7914, 2183, -7875, -2326, 
--7832, 2467, -7789, -2608, 7741, 2746, -7692, -2886, 7639, 3022, -7586, -3159, 7529, 3293, -7471, -3427, 7408, 3559, -7346, -3691, 7279, 3819, -7212, -3949, 7141, 4074, -7070, -4201, 6994, 4324, 
---6919, -4447, 6839, 4567, -6759, -4687, 6676, 4804, -6592, -4921, 6505, 5034, -6417, -5148, 6326, 5257, -6235, -5368, 6140, 5474, -6045, -5580, 5947, 5683, -5849, -5786, 5748, 5885, -5646, -5984, 
--5542, 6079, -5437, -6174, 5330, 6265, -5222, -6356, 5112, 6443, -5002, -6530, 4889, 6613, -4776, -6696, 4660, 6775, -4545, -6854, 4427, 6928, -4310, -7003, 4189, 7073, -4070, -7144, 3947, 7210, 
---3826, -7276, 3701, 7337, -3578, -7399, 3452, 7456, -3327, -7513, 3199, 7566, -3073, -7619, 2944, 7667, -2816, -7716, 2686, 7760, -2557, -7803, 2426, 7843, -2296, -7882, 2163, 7917, -2033, -7952, 
--1899, 7983, -1768, -8013, 1634, 8039, -1502, -8065, 1368, 8086, -1235, -8108, 1101, 8125, -968, -8142, 833, 8155, -701, -8167, 566, 8175, -433, -8183, 299, 8187, -166, -8191, 32, 8190, 
--101, -8190, -234, 8185, 366, -8180, -500, 8171, 631, -8162, -763, 8148, 894, -8135, -1026, 8118, 1155, -8100, -1286, 8078, 1414, -8057, -1544, 8031, 1671, -8005, -1800, 7976, 1926, -7946, 
---2053, 7913, 2178, -7879, -2304, 7841, 2427, -7804, -2551, 7763, 2673, -7722, -2795, 7677, 2915, -7632, -3036, 7583, 3154, -7535, -3273, 7483, 3389, -7431, -3506, 7375, 3620, -7320, -3735, 7260, 
--3847, -7202, -3959, 7139, 4069, -7077, -4179, 7012, 4287, -6947, -4395, 6878, 4500, -6810, -4605, 6738, 4708, -6667, -4811, 6592, 4911, -6518, -5011, 6441, 5108, -6364, -5206, 6284, 5301, -6204, 
---5396, 6121, 5488, -6039, -5580, 5954, 5669, -5869, -5759, 5782, 5845, -5695, -5931, 5605, 6014, -5515, -6098, 5423, 6178, -5332, -6259, 5237, 6336, -5144, -6413, 5048, 6487, -4952, -6562, 4854, 
--6633, -4757, -6704, 4657, 6772, -4558, -6840, 4456, 6905, -4355, -6970, 4252, 7031, -4150, -7093, 4045, 7151, -3942, -7210, 3836, 7264, -3731, -7320, 3623, 7371, -3517, -7423, 3409, 7472, -3302, 
---7520, 3192, 7566, -3084, -7611, 2973, 7653, -2864, -7695, 2753, 7733, -2643, -7772, 2531, 7807, -2421, -7843, 2308, 7875, -2197, -7907, 2084, 7935, -1972, -7964, 1858, 7990, -1747, -8015, 1632, 
--8037, -1520, -8060, 1406, 8079, -1294, -8098, 1179, 8113, -1067, -8129, 952, 8141, -840, -8154, 725, 8163, -613, -8173, 499, 8179, -386, -8185, 272, 8188, -160, -8191, 47, 8190, 65, 
---8191, -178, 8187, 289, -8184, -402, 8178, 513, -8172, -625, 8162, 735, -8153, -847, 8141, 956, -8129, -1067, 8113, 1176, -8098, -1286, 8080, 1394, -8062, -1503, 8041, 1610, -8021, -1718, 
--7997, 1824, -7973, -1931, 7947, 2036, -7921, -2142, 7891, 2246, -7862, -2351, 7830, 2454, -7799, -2558, 7764, 2659, -7730, -2761, 7693, 2861, -7656, -2963, 7617, 3061, -7578, -3161, 7535, 3258, 
---7494, -3357, 7449, 3452, -7406, -3549, 7359, 3643, -7313, -3739, 7264, 3831, -7215, -3925, 7164, 4016, -7113, -4108, 7060, 4197, -7007, -4288, 6952, 4375, -6897, -4464, 6839, 4549, -6783, -4636, 
--6723, 4720, -6664, -4805, 6603, 4888, -6542, -4971, 6479, 5051, -6417, -5132, 6351, 5211, -6287, -5290, 6221, 5366, -6155, -5444, 6086, 5518, -6019, -5594, 5949, 5666, -5880, -5740, 5808, 5810, 
---5738, -5882, 5665, 5950, -5593, -6019, 5518, 6086, -5445, -6153, 5369, 6217, -5295, -6283, 5217, 6345, -5142, -6408, 5063, 6468, -4986, -6529, 4907, 6587, -4829, -6646, 4748, 6702, -4669, -6758, 
--4588, 6812, -4507, -6867, 4425, 6918, -4344, -6971, 4260, 7020, -4179, -7070, 4094, 7118, -4012, -7166, 3926, 7211, -3843, -7257, 3757, 7300, -3673, -7343, 3587, 7384, -3502, -7426, 3415, 7464, 
---3329, -7504, 3242, 7540, -3156, -7577, 3068, 7612, -2981, -7647, 2893, 7679, -2806, -7712, 2717, 7742, -2630, -7773, 2541, 7800, -2454, -7829, 2364, 7855, -2277, -7882, 2187, 7905, -2099, -7930, 
--2009, 7951, -1921, -7974, 1831, 7993, -1743, -8013, 1653, 8031, -1565, -8049, 1475, 8064, -1387, -8081, 1297, 8094, -1209, -8108, 1119, 8120, -1032, -8132, 942, 8141, -854, -8151, 765, 8159, 
---677, -8167, 588, 8172, -500, -8179, 411, 8182, -324, -8187, 236, 8188, -149, -8191, 60, 8190, 26, -8191, -114, 8189, 200, -8188, -287, 8184, 373, -8181, -460, 8175, 545, -8170, 
---631, 8163, 716, -8156, -802, 8147, 886, -8139, -971, 8128, 1055, -8118, -1140, 8105, 1222, -8093, -1306, 8079, 1388, -8066, -1472, 8050, 1553, -8035, -1636, 8017, 1717, -8001, -1799, 7981, 
--1879, -7963, -1960, 7943, 2039, -7923, -2120, 7901, 2198, -7880, -2278, 7856, 2355, -7834, -2434, 7808, 2511, -7784, -2589, 7758, 2665, -7733, -2742, 7705, 2817, -7678, -2893, 7649, 2967, -7621, 
---3042, 7590, 3115, -7561, -3190, 7529, 3262, -7498, -3335, 7465, 3406, -7433, -3478, 7399, 3548, -7366, -3620, 7330, 3689, -7296, -3759, 7259, 3827, -7224, -3897, 7186, 3964, -7150, -4032, 7111, 
--4098, -7073, -4165, 7033, 4230, -6995, -4296, 6954, 4360, -6914, -4425, 6872, 4488, -6832, -4552, 6789, 4613, -6747, -4676, 6703, 4737, -6661, -4799, 6616, 4858, -6573, -4919, 6527, 4977, -6483, 
---5036, 6437, 5093, -6392, -5152, 6345, 5208, -6299, -5265, 6251, 5320, -6205, -5376, 6156, 5430, -6109, -5485, 6059, 5537, -6011, -5591, 5961, 5643, -5913, -5695, 5862, 5745, -5813, -5797, 5762, 
--5846, -5712, -5896, 5660, 5944, -5610, -5994, 5557, 6040, -5506, -6088, 5453, 6134, -5402, -6181, 5349, 6225, -5297, -6271, 5243, 6314, -5191, -6359, 5136, 6401, -5083, -6445, 5029, 6486, -4976, 
---6528, 4920, 6568, -4867, -6609, 4811, 6648, -4758, -6688, 4702, 6726, -4648, -6765, 4591, 6801, -4537, -6839, 4481, 6874, -4426, -6911, 4369, 6945, -4314, -6981, 4257, 7014, -4202, -7048, 4145, 
--7080, -4090, -7114, 4033, 7145, -3977, -7177, 3920, 7207, -3864, -7238, 3806, 7267, -3751, -7297, 3693, 7325, -3637, -7354, 3579, 7381, -3523, -7409, 3466, 7434, -3410, -7461, 3352, 7486, -3296, 
---7512, 3238, 7535, -3182, -7560, 3124, 7583, -3068, -7607, 3010, 7628, -2954, -7651, 2896, 7672, -2840, -7694, 2782, 7714, -2726, -7735, 2668, 7753, -2613, -7773, 2555, 7791, -2499, -7810, 2442, 
--7827, -2386, -7845, 2329, 7861, -2273, -7878, 2216, 7893, -2161, -7909, 2104, 7923, -2048, -7939, 1991, 7952, -1936, -7966, 1880, 7978, -1825, -7992, 1768, 8003, -1714, -8016, 1657, 8027, -1603, 
---8039, 1547, 8048, -1493, -8059, 1437, 8068, -1383, -8079, 1328, 8087, -1274, -8096, 1219, 8103, -1165, -8112, 1110, 8118, -1057, -8127, 1002, 8132, -950, -8139, 895, 8144, -843, -8151, 789, 
--8155, -737, -8161, 683, 8164, -631, -8169, 578, 8172, -526, -8176, 473, 8178, -422, -8182, 369, 8183, -319, -8186, 266, 8187, -216, -8189, 164, 8189, -114, -8191, 62, 8190, -13, 
---8191, -39, 8190, 88, -8191, -139, 8189, 187, -8189, -238, 8186, 286, -8186, -336, 8183, 384, -8181, -434, 8178, 481, -8176, -530, 8172, 577, -8169, -626, 8165, 673, -8162, -721, 
--8157, 767, -8153, -815, 8148, 861, -8144, -909, 8137, 954, -8133, -1001, 8126, 1046, -8121, -1092, 8114, 1137, -8109, -1183, 8101, 1227, -8096, -1272, 8088, 1316, -8081, -1361, 8073, 1404, 
---8066, -1448, 8058, 1491, -8051, -1535, 8041, 1577, -8034, -1621, 8024, 1662, -8016, -1706, 8007, 1747, -7998, -1790, 7988, 1830, -7980, -1873, 7969, 1913, -7960, -1954, 7949, 1994, -7940, -2035, 
--7929, 2074, -7919, -2115, 7907, 2154, -7898, -2194, 7886, 2232, -7876, -2272, 7864, 2310, -7853, -2349, 7841, 2387, -7830, -2426, 7817, 2462, -7807, -2501, 7794, 2537, -7783, -2575, 7769, 2610, 
---7758, -2648, 7745, 2683, -7733, -2720, 7720, 2755, -7708, -2791, 7694, 2825, -7682, -2861, 7668, 2895, -7656, -2931, 7642, 2964, -7630, -2999, 7615, 3032, -7603, -3066, 7588, 3098, -7576, -3132, 
--7561, 3164, -7549, -3198, 7534, 3229, -7521, -3262, 7506, 3293, -7493, -3326, 7478, 3356, -7465, -3388, 7450, 3418, -7437, -3450, 7422, 3479, -7409, -3510, 7393, 3539, -7380, -3570, 7365, 3598, 
---7351, -3629, 7336, 3657, -7323, -3686, 7307, 3714, -7294, -3743, 7278, 3770, -7265, -3799, 7249, 3826, -7236, -3854, 7220, 3880, -7207, -3908, 7191, 3934, -7178, -3961, 7162, 3986, -7148, -4013, 
--7133, 4038, -7119, -4065, 7104, 4089, -7090, -4115, 7075, 4139, -7061, -4165, 7046, 4188, -7032, -4214, 7017, 4237, -7003, -4261, 6988, 4284, -6974, -4308, 6959, 4330, -6946, -4354, 6930, 4376, 
---6917, -4400, 6902, 4421, -6889, -4444, 6873, 4465, -6860, -4488, 6845, 4508, -6832, -4530, 6817, 4550, -6804, -4572, 6789, 4592, -6776, -4613, 6761, 4632, -6749, -4653, 6734, 4672, -6721, -4693, 
--6706, 4711, -6694, -4731, 6679, 4749, -6667, -4769, 6653, 4787, -6640, -4806, 6626, 4823, -6614, -4842, 6600, 4859, -6588, -4878, 6574, 4894, -6562, -4913, 6548, 4929, -6536, -4947, 6522, 4962, 
---6511, -4980, 6497, 4995, -6486, -5012, 6472, 5027, -6461, -5044, 6448, 5058, -6437, -5075, 6424, 5089, -6413, -5105, 6400, 5119, -6389, -5134, 6376, 5148, -6366, -5163, 6353, 5176, -6343, -5191, 
--6330, 5204, -6320, -5218, 6308, 5231, -6298, -5245, 6286, 5257, -6276, -5271, 6264, 5283, -6255, -5296, 6243, 5308, -6234, -5321, 6222, 5332, -6213, -5345, 6202, 5355, -6193, -5368, 6182, 5378, 
---6173, -5390, 6163, 5400, -6154, -5412, 6143, 5422, -6135, -5433, 6125, 5443, -6117, -5454, 6107, 5463, -6099, -5474, 6089, 5482, -6081, -5493, 6072, 5501, -6064, -5512, 6055, 5520, -6048, -5530, 
--6039, 5537, -6032, -5547, 6023, 5554, -6016, -5564, 6008, 5571, -6001, -5580, 5993, 5587, -5987, -5595, 5978, 5602, -5973, -5610, 5965, 5616, -5959, -5624, 5951, 5630, -5946, -5638, 5939, 5644, 
---5933, -5651, 5926, 5657, -5921, -5664, 5914, 5669, -5910, -5676, 5903, 5680, -5899, -5687, 5892, 5691, -5888, -5698, 5882, 5702, -5878, -5708, 5873, 5712, -5869, -5717, 5863, 5721, -5860, -5726, 
--5855, 5729, -5852, -5735, 5847, 5738, -5844, -5742, 5839, 5745, -5837, -5750, 5832, 5752, -5830, -5756, 5826, 5758, -5824, -5762, 5820, 5764, -5818, -5768, 5815, 5769, -5813, -5773, 5810, 5774, 
---5809, -5777, 5806, 5778, -5805, -5781, 5802, 5782, -5801, -5784, 5799, 5785, -5798, -5787, 5796, 5787, -5796, -5789, 5794, 5789, -5794, -5791, 5793, 5790, -5793, -5792, 5792, 5791, -5793, -5792, 
--5791, 5791, -5792, -5792, 5792, 5791, -5793, -5792, 5792, 5790, -5794, -5790, 5794, 5789, -5796, -5789, 5796, 5787, -5798, -5786, 5798, 5784, -5800, -5784, 5801, 5781, -5804, -5780, 5805, 5777, 
---5808, -5776, 5809, 5773, -5812, -5772, 5813, 5768, -5817, -5767, 5819, 5763, -5822, -5761, 5824, 5757, -5828, -5755, 5831, 5750, -5835, -5748, 5837, 5743, -5842, -5740, 5845, 5736, -5850, -5732, 
--5853, 5727, -5858, -5724, 5861, 5718, -5867, -5715, 5870, 5709, -5876, -5705, 5880, 5699, -5886, -5695, 5890, 5689, -5896, -5684, 5900, 5677, -5907, -5673, 5912, 5666, -5918, -5661, 5923, 5653, 
---5930, -5648, 5935, 5640, -5943, -5635, 5948, 5627, -5956, -5621, 5961, 5613, -5969, -5607, 5975, 5598, -5983, -5591, 5989, 5583, -5997, -5576, 6004, 5567, -6012, -5560, 6019, 5550, -6028, -5543, 
--6035, 5533, -6044, -5525, 6051, 5515, -6060, -5507, 6068, 5497, -6077, -5488, 6085, 5478, -6094, -5469, 6102, 5458, -6112, -5449, 6120, 5438, -6130, -5428, 6139, 5417, -6149, -5407, 6158, 5395, 
---6168, -5385, 6177, 5372, -6188, -5362, 6197, 5349, -6208, -5339, 6217, 5326, -6228, -5315, 6238, 5301, -6249, -5290, 6259, 5276, -6271, -5265, 6280, 5251, -6292, -5238, 6302, 5224, -6314, -5212, 
--6325, 5197, -6337, -5184, 6347, 5169, -6360, -5156, 6370, 5141, -6383, -5127, 6394, 5111, -6407, -5097, 6418, 5081, -6431, -5067, 6442, 5051, -6455, -5036, 6466, 5019, -6479, -5004, 6491, 4987, 
---6504, -4971, 6516, 4954, -6530, -4938, 6541, 4920, -6555, -4904, 6567, 4886, -6581, -4869, 6593, 4850, -6607, -4833, 6619, 4814, -6634, -4797, 6646, 4778, -6660, -4760, 6673, 4740, -6687, -4722, 
--6700, 4701, -6714, -4683, 6727, 4662, -6742, -4643, 6754, 4622, -6769, -4603, 6782, 4581, -6797, -4562, 6810, 4540, -6825, -4520, 6838, 4497, -6853, -4477, 6866, 4454, -6881, -4433, 6895, 4410, 
---6910, -4388, 6923, 4365, -6939, -4343, 6952, 4319, -6967, -4297, 6981, 4272, -6996, -4249, 7009, 4225, -7025, -4201, 7038, 4176, -7054, -4153, 7067, 4127, -7083, -4103, 7096, 4076, -7112, -4052, 
--7126, 4025, -7141, -4000, 7155, 3973, -7170, -3948, 7184, 3920, -7199, -3895, 7213, 3867, -7228, -3840, 7242, 3812, -7257, -3785, 7271, 3756, -7286, -3729, 7300, 3700, -7315, -3672, 7329, 3642, 
---7344, -3614, 7358, 3584, -7373, -3555, 7386, 3524, -7401, -3495, 7415, 3464, -7430, -3434, 7443, 3403, -7458, -3373, 7471, 3340, -7486, -3310, 7499, 3277, -7514, -3246, 7527, 3213, -7542, -3182, 
--7554, 3148, -7569, -3116, 7582, 3082, -7596, -3049, 7609, 3015, -7623, -2982, 7635, 2947, -7649, -2913, 7662, 2878, -7676, -2844, 7688, 2808, -7701, -2773, 7713, 2737, -7727, -2702, 7738, 2665, 
---7752, -2630, 7763, 2592, -7776, -2556, 7788, 2518, -7801, -2482, 7812, 2443, -7824, -2407, 7835, 2368, -7847, -2330, 7858, 2291, -7870, -2253, 7880, 2213, -7892, -2175, 7902, 2134, -7914, -2095, 
--7923, 2054, -7935, -2015, 7944, 1974, -7955, -1934, 7964, 1892, -7975, -1852, 7983, 1809, -7994, -1769, 8002, 1726, -8012, -1685, 8020, 1641, -8030, -1600, 8037, 1556, -8046, -1514, 8054, 1469, 
---8063, -1427, 8069, 1382, -8078, -1339, 8084, 1293, -8092, -1250, 8098, 1204, -8106, -1160, 8111, 1114, -8118, -1069, 8123, 1023, -8130, -978, 8135, 931, -8141, -885, 8145, 838, -8151, -792, 
--8154, 744, -8160, -698, 8163, 649, -8168, -602, 8170, 553, -8174, -506, 8176, 457, -8180, -409, 8181, 360, -8185, -312, 8185, 261, -8188, -213, 8188, 162, -8190, -114, 8190, 63, 
---8191, -13, 8190, -38, -8191, 88, 8190, -139, -8190, 189, 8188, -242, -8187, 292, 8184, -344, -8183, 395, 8180, -448, -8178, 499, 8174, -552, -8171, 604, 8166, -657, -8163, 709, 
--8157, -763, -8153, 815, 8147, -870, -8142, 922, 8135, -977, -8130, 1029, 8122, -1084, -8116, 1137, 8107, -1192, -8100, 1246, 8091, -1301, -8083, 1355, 8073, -1411, -8064, 1464, 8053, -1520, 
---8044, 1575, 8032, -1631, -8022, 1685, 8009, -1742, -7998, 1796, 7985, -1853, -7973, 1908, 7958, -1964, -7946, 2019, 7930, -2076, -7917, 2132, 7901, -2189, -7886, 2244, 7869, -2301, -7853, 2357, 
--7835, -2414, -7819, 2470, 7800, -2528, -7783, 2583, 7763, -2641, -7744, 2697, 7724, -2755, -7704, 2811, 7683, -2868, -7662, 2924, 7640, -2982, -7618, 3038, 7595, -3096, -7572, 3152, 7548, -3210, 
---7524, 3266, 7498, -3324, -7474, 3380, 7447, -3438, -7422, 3494, 7394, -3552, -7368, 3608, 7339, -3666, -7312, 3721, 7282, -3779, -7253, 3835, 7222, -3892, -7193, 3948, 7160, -4005, -7130, 4061, 
--7097, -4118, -7065, 4173, 7031, -4230, -6998, 4285, 6962, -4342, -6929, 4397, 6892, -4454, -6857, 4508, 6819, -4565, -6783, 4619, 6745, -4675, -6707, 4729, 6668, -4785, -6629, 4839, 6588, -4894, 
---6549, 4947, 6507, -5003, -6466, 5056, 6423, -5110, -6381, 5163, 6336, -5217, -6293, 5269, 6248, -5323, -6204, 5375, 6157, -5428, -6112, 5479, 6064, -5532, -6018, 5583, 5969, -5635, -5921, 5685, 
--5871, -5737, -5822, 5787, 5771, -5838, -5721, 5887, 5668, -5938, -5617, 5986, 5564, -6036, -5512, 6083, 5457, -6133, -5404, 6180, 5348, -6228, -5293, 6274, 5236, -6322, -5180, 6368, 5122, -6415, 
---5066, 6460, 5006, -6506, -4948, 6550, 4888, -6595, -4829, 6638, 4767, -6683, -4707, 6725, 4644, -6768, -4583, 6810, 4519, -6852, -4457, 6893, 4392, -6934, -4329, 6974, 4263, -7014, -4198, 7053, 
--4131, -7092, -4066, 7130, 3997, -7168, -3931, 7204, 3862, -7242, -3794, 7277, 3724, -7314, -3655, 7347, 3584, -7383, -3514, 7415, 3442, -7450, -3371, 7481, 3298, -7514, -3226, 7544, 3152, -7576, 
---3079, 7605, 3004, -7635, -2930, 7663, 2854, -7692, -2780, 7718, 2703, -7746, -2627, 7771, 2549, -7797, -2473, 7821, 2394, -7845, -2317, 7868, 2238, -7891, -2159, 7912, 2079, -7933, -2000, 7953, 
--1919, -7973, -1839, 7991, 1757, -8009, -1677, 8026, 1594, -8043, -1513, 8057, 1430, -8073, -1348, 8086, 1264, -8100, -1181, 8111, 1097, -8123, -1014, 8133, 928, -8143, -844, 8151, 758, -8160, 
---674, 8166, 588, -8173, -503, 8178, 416, -8183, -331, 8185, 243, -8189, -157, 8190, 69, -8191, 17, 8190, -105, -8190, 192, 8187, -280, -8185, 367, 8180, -456, -8176, 543, 8169, 
---633, -8164, 720, 8155, -810, -8147, 897, 8136, -987, -8126, 1075, 8114, -1165, -8102, 1253, 8087, -1343, -8073, 1431, 8056, -1521, -8041, 1609, 8022, -1699, -8004, 1787, 7983, -1877, -7963, 
--1965, 7940, -2055, -7918, 2143, 7893, -2232, -7869, 2320, 7842, -2409, -7816, 2497, 7786, -2586, -7758, 2673, 7726, -2762, -7696, 2849, 7662, -2938, -7630, 3024, 7594, -3112, -7559, 3198, 7521, 
---3286, -7485, 3372, 7445, -3459, -7405, 3544, 7363, -3630, -7322, 3715, 7278, -3801, -7234, 3884, 7188, -3970, -7142, 4052, 7094, -4137, -7046, 4219, 6995, -4303, -6945, 4384, 6892, -4467, -6840, 
--4547, 6785, -4629, -6731, 4708, 6673, -4789, -6617, 4867, 6558, -4947, -6499, 5024, 6438, -5103, -6377, 5179, 6313, -5257, -6251, 5331, 6185, -5408, -6120, 5481, 6052, -5556, -5985, 5628, 5915, 
---5702, -5847, 5773, 5775, -5845, -5704, 5914, 5630, -5984, -5557, 6052, 5481, -6121, -5406, 6187, 5328, -6255, -5251, 6319, 5171, -6385, -5092, 6447, 5010, -6511, -4930, 6572, 4846, -6634, -4763, 
--6693, 4678, -6753, -4594, 6811, 4506, -6869, -4420, 6924, 4331, -6980, -4243, 7033, 4152, -7087, -4062, 7138, 3970, -7190, -3879, 7239, 3784, -7289, -3691, 7335, 3596, -7383, -3501, 7427, 3404, 
---7472, -3308, 7514, 3209, -7557, -3112, 7597, 3011, -7637, -2913, 7674, 2811, -7712, -2711, 7747, 2608, -7782, -2506, 7814, 2402, -7847, -2299, 7876, 2194, -7906, -2090, 7933, 1983, -7961, -1878, 
--7985, 1771, -8009, -1665, 8031, 1556, -8053, -1449, 8071, 1339, -8090, -1232, 8106, 1121, -8122, -1012, 8134, 901, -8148, -792, 8157, 680, -8168, -570, 8174, 457, -8182, -346, 8185, 233, 
---8190, -122, 8190, 9, -8191, 103, 8189, -217, -8187, 329, 8181, -443, -8176, 555, 8168, -670, -8159, 782, 8147, -896, -8136, 1009, 8121, -1123, -8106, 1236, 8088, -1350, -8070, 1463, 
--8048, -1577, -8027, 1689, 8002, -1803, -7978, 1915, 7950, -2028, -7922, 2140, 7891, -2253, -7859, 2364, 7825, -2476, -7790, 2587, 7752, -2699, -7715, 2808, 7674, -2919, -7633, 3028, 7588, -3139, 
---7544, 3246, 7496, -3356, -7448, 3463, 7397, -3571, -7346, 3677, 7292, -3784, -7238, 3888, 7180, -3994, -7123, 4097, 7062, -4202, -7001, 4303, 6937, -4406, -6873, 4506, 6806, -4608, -6739, 4706, 
--6668, -4806, -6598, 4903, 6524, -5000, -6451, 5095, 6374, -5191, -6298, 5284, 6218, -5378, -6139, 5469, 6056, -5561, -5973, 5649, 5888, -5739, -5802, 5825, 5713, -5912, -5625, 5996, 5534, -6081, 
---5443, 6162, 5348, -6245, -5254, 6323, 5157, -6403, -5060, 6479, 4961, -6556, -4861, 6629, 4759, -6703, -4657, 6774, 4552, -6845, -4448, 6912, 4340, -6980, -4234, 7044, 4124, -7109, -4015, 7170, 
--3903, -7232, -3791, 7290, 3677, -7348, -3564, 7402, 3447, -7457, -3332, 7508, 3213, -7560, -3096, 7607, 2975, -7655, -2856, 7699, 2734, -7743, -2613, 7783, 2489, -7824, -2366, 7860, 2241, -7896, 
---2116, 7929, 1989, -7962, -1864, 7990, 1735, -8019, -1608, 8044, 1479, -8068, -1351, 8089, 1220, -8110, -1091, 8126, 959, -8143, -829, 8155, 697, -8167, -566, 8175, 432, -8183, -301, 8187, 
--167, -8191, -35, 8190, -99, -8190, 232, 8185, -366, -8180, 499, 8171, -634, -8162, 767, 8148, -901, -8134, 1034, 8116, -1169, -8098, 1301, 8075, -1435, -8053, 1568, 8026, -1702, -7999, 
--1833, 7967, -1966, -7935, 2097, 7900, -2230, -7863, 2360, 7823, -2492, -7782, 2621, 7737, -2752, -7692, 2880, 7643, -3009, -7593, 3136, 7540, -3264, -7486, 3389, 7427, -3516, -7369, 3639, 7306, 
---3764, -7243, 3886, 7176, -4009, -7109, 4129, 7038, -4250, -6966, 4368, 6891, -4487, -6815, 4602, 6735, -4719, -6655, 4832, 6571, -4946, -6487, 5056, 6399, -5168, -6311, 5276, 6219, -5384, -6127, 
--5489, 6031, -5595, -5935, 5697, 5835, -5799, -5735, 5898, 5631, -5997, -5528, 6092, 5420, -6188, -5313, 6280, 5202, -6372, -5092, 6461, 4977, -6549, -4863, 6634, 4745, -6718, -4628, 6799, 4507, 
---6880, -4386, 6956, 4262, -7033, -4138, 7105, 4011, -7177, -3885, 7245, 3755, -7313, -3625, 7377, 3493, -7440, -3361, 7499, 3225, -7558, -3091, 7613, 2953, -7667, -2817, 7716, 2677, -7765, -2538, 
--7810, 2396, -7854, -2255, 7894, 2111, -7933, -1969, 7968, 1823, -8002, -1679, 8032, 1532, -8061, -1386, 8085, 1238, -8108, -1091, 8127, 941, -8145, -793, 8159, 642, -8172, -493, 8180, 342, 
---8187, -192, 8190, 41, -8191, 110, 8188, -262, -8185, 412, 8176, -565, -8166, 715, 8152, -867, -8137, 1018, 8117, -1170, -8096, 1320, 8071, -1471, -8044, 1621, 8013, -1772, -7981, 1920, 
--7944, -2070, -7906, 2218, 7863, -2367, -7820, 2513, 7771, -2660, -7722, 2805, 7668, -2951, -7613, 3094, 7554, -3239, -7493, 3380, 7428, -3522, -7362, 3661, 7291, -3801, -7220, 3938, 7144, -4075, 
---7067, 4209, 6985, -4344, -6903, 4475, 6816, -4607, -6729, 4735, 6637, -4864, -6544, 4989, 6447, -5115, -6349, 5236, 6247, -5358, -6144, 5476, 6037, -5594, -5930, 5708, 5818, -5822, -5706, 5932, 
--5589, -6042, -5472, 6148, 5351, -6253, -5230, 6355, 5105, -6456, -4979, 6552, 4850, -6648, -4720, 6740, 4587, -6831, -4453, 6918, 4316, -7004, -4179, 7086, 4038, -7167, -3897, 7243, 3752, -7318, 
---3608, 7389, 3460, -7458, -3313, 7523, 3162, -7587, -3012, 7646, 2859, -7704, -2706, 7758, 2550, -7810, -2394, 7857, 2236, -7902, -2078, 7943, 1917, -7983, -1758, 8017, 1595, -8050, -1434, 8078, 
--1270, -8105, -1107, 8126, 942, -8146, -777, 8161, 611, -8174, -446, 8182, 278, -8189, -113, 8190, -55, -8190, 221, 8185, -390, -8178, 556, 8165, -724, -8152, 890, 8132, -1058, -8112, 
--1224, 8085, -1391, -8058, 1556, 8025, -1723, -7990, 1887, 7950, -2052, -7909, 2215, 7862, -2379, -7813, 2540, 7760, -2702, -7705, 2861, 7644, -3022, -7582, 3179, 7515, -3336, -7446, 3491, 7372, 
---3646, -7297, 3798, 7216, -3950, -7134, 4099, 7047, -4248, -6959, 4393, 6866, -4539, -6771, 4681, 6671, -4823, -6570, 4960, 6465, -5098, -6358, 5232, 6246, -5365, -6133, 5494, 6015, -5623, -5897, 
--5748, 5773, -5872, -5649, 5991, 5520, -6110, -5391, 6224, 5257, -6338, -5122, 6446, 4983, -6554, -4843, 6657, 4699, -6759, -4555, 6856, 4406, -6952, -4258, 7043, 4105, -7133, -3951, 7217, 3794, 
---7300, -3637, 7378, 3476, -7454, -3316, 7525, 3151, -7595, -2987, 7659, 2819, -7721, -2652, 7778, 2481, -7833, -2311, 7883, 2138, -7930, -1965, 7972, 1790, -8013, -1615, 8047, 1437, -8080, -1261, 
--8106, 1081, -8131, -903, 8150, 722, -8167, -543, 8178, 361, -8187, -181, 8190, -1, -8191, 182, 8186, -365, -8179, 546, 8166, -728, -8150, 909, 8129, -1091, -8106, 1271, 8076, -1453, 
---8045, 1631, 8008, -1812, -7968, 1989, 7922, -2168, -7875, 2344, 7821, -2521, -7765, 2695, 7703, -2870, -7640, 3041, 7570, -3213, -7499, 3381, 7421, -3550, -7342, 3716, 7256, -3881, -7169, 4043, 
--7076, -4205, -6982, 4363, 6881, -4521, -6779, 4674, 6672, -4828, -6563, 4976, 6448, -5125, -6331, 5269, 6210, -5412, -6087, 5551, 5958, -5689, -5828, 5822, 5693, -5954, -5557, 6081, 5416, -6207, 
---5274, 6328, 5127, -6447, -4979, 6561, 4826, -6674, -4672, 6782, 4514, -6887, -4355, 6987, 4191, -7086, -4027, 7179, 3859, -7270, -3691, 7355, 3518, -7438, -3345, 7515, 3168, -7590, -2991, 7659, 
--2811, -7726, -2631, 7787, 2447, -7846, -2263, 7898, 2076, -7948, -1890, 7991, 1701, -8032, -1512, 8067, 1320, -8099, -1130, 8125, 936, -8148, -744, 8165, 549, -8179, -356, 8186, 160, -8191, 
--34, 8189, -230, -8185, 424, 8174, -620, -8160, 814, 8140, -1010, -8116, 1203, 8087, -1398, -8054, 1590, 8015, -1784, -7973, 1974, 7925, -2166, -7873, 2355, 7816, -2544, -7755, 2730, 7688, 
---2917, -7619, 3100, 7543, -3284, -7464, 3464, 7379, -3644, -7292, 3820, 7198, -3996, -7102, 4168, 6999, -4339, -6895, 4506, 6784, -4673, -6671, 4835, 6551, -4996, -6430, 5152, 6303, -5308, -6174, 
--5458, 6039, -5607, -5902, 5751, 5760, -5894, -5616, 6031, 5466, -6167, -5315, 6297, 5159, -6426, -5001, 6548, 4838, -6669, -4674, 6784, 4505, -6896, -4335, 7003, 4160, -7107, -3985, 7205, 3804, 
---7301, -3624, 7390, 3438, -7477, -3253, 7557, 3063, -7635, -2873, 7705, 2680, -7774, -2486, 7835, 2289, -7893, -2092, 7945, 1891, -7993, -1691, 8035, 1488, -8073, -1286, 8105, 1080, -8133, -876, 
--8154, 669, -8172, -464, 8183, 255, -8190, -49, 8190, -160, -8187, 366, 8177, -575, -8163, 782, 8142, -990, -8118, 1196, 8087, -1403, -8052, 1607, 8010, -1813, -7965, 2016, 7912, -2219, 
---7856, 2419, 7793, -2620, -7727, 2818, 7654, -3015, -7577, 3209, 7494, -3403, -7407, 3593, 7313, -3782, -7217, 3968, 7113, -4152, -7007, 4333, 6894, -4512, -6778, 4687, 6656, -4860, -6531, 5029, 
--6399, -5196, -6265, 5358, 6124, -5518, -5982, 5673, 5833, -5826, -5682, 5973, 5525, -6119, -5366, 6258, 5201, -6395, -5035, 6526, 4863, -6655, -4689, 6777, 4510, -6896, -4330, 7009, 4145, -7119, 
---3958, 7222, 3767, -7323, -3575, 7416, 3378, -7506, -3181, 7589, 2979, -7669, -2777, 7742, 2571, -7811, -2365, 7873, 2155, -7931, -1945, 7981, 1732, -8029, -1519, 8068, 1303, -8104, -1088, 8132, 
--870, -8156, -653, 8172, 434, -8185, -216, 8190, -5, -8191, 223, 8184, -444, -8173, 662, 8154, -883, -8131, 1100, 8101, -1320, -8066, 1536, 8024, -1753, -7977, 1968, 7923, -2183, -7865, 
--2395, 7799, -2607, -7730, 2815, 7652, -3024, -7571, 3228, 7483, -3433, -7390, 3633, 7291, -3832, -7187, 4027, 7076, -4221, -6962, 4410, 6841, -4598, -6716, 4780, 6585, -4961, -6450, 5137, 6308, 
---5311, -6163, 5479, 6012, -5645, -5858, 5805, 5697, -5963, -5534, 6114, 5365, -6263, -5193, 6405, 5015, -6545, -4836, 6677, 4650, -6807, -4463, 6929, 4270, -7049, -4076, 7161, 3876, -7269, -3675, 
--7370, 3469, -7468, -3263, 7557, 3051, -7643, -2840, 7722, 2623, -7796, -2407, 7862, 2186, -7924, -1966, 7978, 1741, -8028, -1518, 8069, 1291, -8106, -1064, 8135, 835, -8160, -607, 8176, 376, 
---8187, -146, 8190, -85, -8189, 315, 8179, -547, -8165, 777, 8142, -1008, -8114, 1236, 8078, -1466, -8038, 1693, 7989, -1920, -7935, 2145, 7873, -2369, -7807, 2590, 7732, -2811, -7653, 3028, 
--7566, -3245, -7474, 3457, 7375, -3669, -7271, 3876, 7159, -4081, -7043, 4282, 6920, -4481, -6792, 4675, 6657, -4867, -6518, 5053, 6372, -5237, -6223, 5415, 6066, -5591, -5906, 5760, 5739, -5927, 
---5569, 6087, 5392, -6243, -5212, 6393, 5027, -6540, -4838, 6679, 4644, -6814, -4447, 6942, 4245, -7067, -4040, 7183, 3831, -7295, -3619, 7400, 3403, -7500, -3185, 7592, 2963, -7679, -2740, 7758, 
--2512, -7833, -2284, 7898, 2052, -7959, -1820, 8012, 1584, -8059, -1348, 8098, 1110, -8131, -872, 8156, 631, -8176, -391, 8186, 149, -8191, 91, 8188, -334, -8179, 574, 8161, -817, -8138, 
--1056, 8106, -1297, -8068, 1535, 8022, -1774, -7970, 2009, 7909, -2245, -7844, 2477, 7769, -2710, -7689, 2937, 7601, -3165, -7508, 3388, 7406, -3610, -7299, 3827, 7183, -4042, -7064, 4253, 6935, 
---4461, -6803, 4664, 6662, -4865, -6517, 5059, 6364, -5252, -6207, 5437, 6043, -5620, -5875, 5796, 5699, -5968, -5520, 6134, 5334, -6296, -5145, 6450, 4949, -6601, -4751, 6744, 4546, -6882, -4338, 
--7013, 4125, -7139, -3909, 7256, 3688, -7369, -3465, 7474, 3237, -7573, -3007, 7664, 2773, -7749, -2538, 7825, 2298, -7897, -2058, 7958, 1814, -8015, -1570, 8062, 1322, -8103, -1075, 8135, 825, 
---8162, -575, 8178, 323, -8189, -73, 8190, -180, -8186, 431, 8172, -684, -8151, 934, 8122, -1185, -8086, 1434, 8041, -1683, -7990, 1929, 7929, -2175, -7863, 2418, 7787, -2660, -7706, 2898, 
--7615, -3135, -7518, 3368, 7413, -3599, -7302, 3825, 7182, -4050, -7057, 4269, 6923, -4486, -6784, 4696, 6636, -4904, -6484, 5106, 6323, -5305, -6158, 5496, 5985, -5685, -5808, 5866, 5623, -6043, 
---5435, 6213, 5238, -6379, -5039, 6536, 4832, -6689, -4623, 6834, 4407, -6973, -4188, 7104, 3963, -7231, -3735, 7348, 3502, -7459, -3267, 7562, 3027, -7658, -2786, 7746, 2539, -7827, -2292, 7899, 
--2040, -7965, -1788, 8020, 1532, -8070, -1276, 8110, 1017, -8143, -759, 8166, 497, -8183, -237, 8190, -25, -8190, 286, 8180, -549, -8163, 809, 8136, -1071, -8103, 1329, 8059, -1589, -8010, 
--1845, 7949, -2101, -7883, 2354, 7806, -2606, -7723, 2854, 7630, -3100, -7531, 3342, 7422, -3583, -7308, 3818, 7183, -4051, -7053, 4278, 6914, -4503, -6769, 4721, 6615, -4937, -6456, 5145, 6288, 
---5350, -6116, 5548, 5934, -5742, -5748, 5928, 5555, -6110, -5357, 6283, 5151, -6452, -4941, 6612, 4724, -6768, -4504, 6914, 4277, -7055, -4048, 7186, 3811, -7312, -3573, 7428, 3328, -7538, -3082, 
--7638, 2830, -7732, -2577, 7816, 2319, -7893, -2060, 7960, 1797, -8020, -1534, 8070, 1267, -8113, -1000, 8145, 730, -8170, -461, 8184, 189, -8191, 81, 8188, -353, -8177, 623, 8155, -895, 
---8127, 1164, 8087, -1433, -8040, 1700, 7983, -1966, -7918, 2229, 7843, -2491, -7761, 2749, 7668, -3006, -7569, 3257, 7459, -3508, -7343, 3752, 7216, -3995, -7084, 4231, 6941, -4464, -6792, 4691, 
--6634, -4915, -6470, 5131, 6297, -5344, -6118, 5548, 5930, -5749, -5738, 5941, 5537, -6129, -5331, 6308, 5117, -6481, -4899, 6646, 4674, -6805, -4445, 6954, 4208, -7098, -3969, 7231, 3723, -7358, 
---3475, 7475, 3220, -7585, -2963, 7685, 2701, -7778, -2438, 7860, 2169, -7935, -1900, 7998, 1627, -8055, -1353, 8100, 1076, -8138, -799, 8164, 519, -8183, -240, 8190, -41, -8190, 321, 8177, 
---602, -8158, 881, 8127, -1161, -8088, 1437, 8037, -1714, -7980, 1988, 7910, -2261, -7833, 2530, 7745, -2798, -7650, 3060, 7543, -3322, -7429, 3577, 7305, -3831, -7173, 4078, 7031, -4322, -6883, 
--4559, 6724, -4793, -6559, 5020, 6384, -5242, -6203, 5457, 6012, -5667, -5816, 5868, 5611, -6064, -5401, 6251, 5182, -6433, -4959, 6605, 4728, -6771, -4492, 6926, 4249, -7076, -4003, 7215, 3750, 
---7347, -3493, 7468, 3231, -7583, -2966, 7686, 2696, -7781, -2423, 7865, 2146, -7942, -1868, 8006, 1585, -8063, -1303, 8108, 1016, -8145, -730, 8170, 441, -8186, -153, 8190, -137, -8187, 425, 
--8171, -715, -8146, 1003, 8110, -1291, -8065, 1575, 8008, -1860, -7943, 2141, 7866, -2422, -7781, 2697, 7684, -2971, -7580, 3240, 7463, -3507, -7340, 3767, 7204, -4025, -7062, 4276, 6908, -4524, 
---6748, 4764, 6576, -5000, -6399, 5228, 6211, -5451, -6016, 5665, 5812, -5875, -5603, 6075, 5384, -6269, -5160, 6453, 4927, -6631, -4689, 6799, 4444, -6960, -4194, 7110, 3937, -7253, -3677, 7384, 
--3409, -7508, -3139, 7621, 2863, -7725, -2585, 7818, 2301, -7902, -2016, 7974, 1726, -8037, -1436, 8088, 1142, -8131, -848, 8161, 550, -8182, -254, 8190, -45, -8189, 342, 8176, -640, -8153, 
--936, 8118, -1233, -8074, 1527, 8018, -1821, -7952, 2110, 7874, -2399, -7787, 2683, 7688, -2965, -7581, 3242, 7461, -3516, -7333, 3784, 7193, -4049, -7046, 4307, 6886, -4561, -6720, 4807, 6542, 
---5049, -6357, 5282, 6162, -5510, -5960, 5728, 5747, -5941, -5529, 6144, 5301, -6341, -5068, 6527, 4825, -6707, -4578, 6875, 4323, -7037, -4063, 7186, 3796, -7328, -3525, 7458, 3247, -7579, -2967, 
--7688, 2680, -7789, -2391, 7877, 2097, -7956, -1802, 8022, 1502, -8079, -1202, 8123, 898, -8157, -594, 8179, 287, -8190, 18, 8189, -325, -8178, 630, 8153, -937, -8119, 1240, 8071, -1544, 
---8014, 1843, 7944, -2143, -7865, 2437, 7772, -2730, -7671, 3018, 7556, -3303, -7433, 3582, 7297, -3858, -7152, 4127, 6995, -4392, -6830, 4649, 6654, -4902, -6470, 5145, 6274, -5384, -6071, 5613, 
--5858, -5835, -5637, 6048, 5407, -6254, -5171, 6450, 4925, -6638, -4674, 6814, 4413, -6983, -4149, 7140, 3876, -7289, -3599, 7425, 3315, -7552, -3028, 7667, 2735, -7772, -2439, 7864, 2137, -7947, 
---1835, 8016, 1527, -8076, -1219, 8121, 907, -8157, -595, 8179, 280, -8191, 33, 8188, -349, -8176, 662, 8149, -976, -8113, 1287, 8062, -1599, -8002, 1906, 7927, -2213, -7843, 2514, 7745, 
---2814, -7637, 3108, 7516, -3400, -7386, 3684, 7242, -3965, -7090, 4239, 6925, -4508, -6751, 4769, 6565, -5025, -6371, 5271, 6165, -5511, -5952, 5742, 5728, -5965, -5497, 6178, 5256, -6384, -5008, 
--6578, 4751, -6764, -4488, 6938, 4216, -7104, -3940, 7257, 3655, -7400, -3367, 7531, 3071, -7652, -2773, 7760, 2468, -7858, -2161, 7941, 1849, -8015, -1535, 8074, 1217, -8123, -899, 8157, 578, 
---8181, -257, 8190, -67, -8188, 388, 8172, -711, -8145, 1031, 8103, -1352, -8051, 1669, 7984, -1985, -7907, 2296, 7815, -2607, -7713, 2911, 7597, -3213, -7470, 3508, 7330, -3799, -7181, 4083, 
--7018, -4363, -6845, 4633, 6660, -4899, -6467, 5155, 6261, -5405, -6046, 5645, 5821, -5878, -5587, 6100, 5343, -6314, -5092, 6516, 4831, -6710, -4564, 6891, 4288, -7064, -4006, 7223, 3716, -7373, 
---3422, 7509, 3120, -7635, -2815, 7747, 2503, -7848, -2189, 7935, 1870, -8011, -1549, 8072, 1223, -8123, -897, 8158, 568, -8182, -239, 8190, -92, -8187, 421, 8169, -752, -8140, 1079, 8096, 
---1407, -8040, 1731, 7969, -2055, -7887, 2373, 7789, -2689, -7682, 3000, 7559, -3307, -7426, 3607, 7278, -3904, -7121, 4192, 6950, -4476, -6769, 4750, 6574, -5018, -6371, 5277, 6155, -5528, -5931, 
--5769, 5695, -6002, -5451, 6224, 5196, -6437, -4934, 6638, 4662, -6829, -4383, 7008, 4095, -7176, -3803, 7331, 3501, -7475, -3196, 7605, 2883, -7725, -2567, 7829, 2244, -7922, -1920, 8000, 1590, 
---8067, -1259, 8117, 924, -8156, -589, 8180, 251, -8191, 86, 8187, -424, -8170, 761, 8138, -1098, -8093, 1431, 8033, -1764, -7961, 2093, 7874, -2420, -7774, 2741, 7660, -3059, -7534, 3371, 
--7393, -3678, -7241, 3978, 7075, -4273, -6899, 4559, 6708, -4839, -6508, 5109, 6294, -5372, -6071, 5624, 5836, -5868, -5592, 6100, 5337, -6324, -5074, 6535, 4800, -6736, -4519, 6924, 4229, -7102, 
---3932, 7266, 3627, -7419, -3317, 7557, 3000, -7684, -2678, 7795, 2350, -7895, -2020, 7978, 1684, -8050, -1346, 8106, 1004, -8149, -662, 8176, 317, -8190, 27, 8188, -373, -8173, 717, 8142, 
---1062, -8098, 1403, 8038, -1743, -7965, 2079, 7876, -2413, -7775, 2741, 7658, -3067, -7529, 3385, 7385, -3699, -7229, 4005, 7058, -4305, -6876, 4596, 6680, -4881, -6474, 5155, 6253, -5422, -6024, 
--5678, 5781, -5925, -5529, 6159, 5266, -6385, -4994, 6597, 4712, -6799, -4423, 6987, 4123, -7164, -3818, 7327, 3503, -7477, -3184, 7613, 2857, -7736, -2527, 7843, 2190, -7938, -1850, 8017, 1505, 
---8082, -1159, 8131, 809, -8167, -459, 8186, 106, -8191, 246, 8180, -599, -8155, 949, 8113, -1300, -8058, 1647, 7986, -1992, -7901, 2332, 7799, -2670, -7685, 3002, 7554, -3329, -7411, 3649, 
--7252, -3964, -7081, 4270, 6895, -4570, -6698, 4859, 6486, -5142, -6264, 5413, 6028, -5676, -5782, 5926, 5524, -6167, -5256, 6395, 4977, -6613, -4690, 6816, 4392, -7008, -4087, 7186, 3773, -7351, 
---3453, 7501, 3124, -7638, -2792, 7759, 2451, -7868, -2108, 7959, 1759, -8037, -1408, 8098, 1052, -8145, -696, 8174, 336, -8190, 22, 8188, -383, -8172, 741, 8139, -1099, -8091, 1454, 8026, 
---1809, -7948, 2158, 7852, -2505, -7742, 2845, 7616, -3182, -7476, 3511, 7320, -3835, -7152, 4150, 6968, -4459, -6772, 4757, 6560, -5049, -6338, 5328, 6101, -5599, -5854, 5858, 5593, -6107, -5323, 
--6342, 5040, -6567, -4750, 6777, 4448, -6976, -4139, 7159, 3819, -7330, -3494, 7484, 3160, -7626, -2821, 7750, 2475, -7862, -2125, 7956, 1769, -8036, -1411, 8098, 1048, -8145, -685, 8175, 319, 
---8190, 47, 8187, -414, -8170, 779, 8134, -1145, -8084, 1506, 8015, -1867, -7932, 2222, 7831, -2574, -7717, 2920, 7585, -3262, -7439, 3596, 7276, -3924, -7100, 4243, 6908, -4555, -6704, 4857, 
--6484, -5150, -6253, 5431, 6006, -5703, -5750, 5962, 5479, -6211, -5200, 6445, 4907, -6668, -4606, 6875, 4294, -7071, -3975, 7250, 3645, -7416, -3309, 7566, 2965, -7701, -2616, 7819, 2260, -7923, 
---1901, 8008, 1536, -8079, -1169, 8131, 798, -8169, -427, 8187, 53, -8190, 319, 8175, -693, -8144, 1064, 8095, -1435, -8030, 1801, 7947, -2165, -7849, 2523, 7732, -2878, -7602, 3225, 7453, 
---3568, -7290, 3901, 7110, -4228, -6918, 4544, 6708, -4853, -6486, 5150, 6248, -5438, -5999, 5713, 5736, -5978, -5462, 6228, 5174, -6468, -4877, 6691, 4567, -6903, -4250, 7098, 3922, -7280, -3587, 
--7445, 3242, -7595, -2892, 7728, 2533, -7846, -2171, 7946, 1803, -8030, -1432, 8095, 1056, -8145, -679, 8176, 299, -8191, 80, 8186, -461, -8166, 839, 8126, -1218, -8070, 1592, 7995, -1965, 
---7904, 2332, 7795, -2696, -7670, 3053, 7527, -3405, -7369, 3747, 7193, -4084, -7004, 4410, 6797, -4729, -6577, 5035, 6340, -5332, -6092, 5616, 5828, -5890, -5553, 6149, 5264, -6397, -4965, 6629, 
--4654, -6848, -4333, 7051, 4001, -7239, -3662, 7410, 3313, -7567, -2958, 7705, 2595, -7828, -2227, 7932, 1853, -8021, -1476, 8089, 1094, -8142, -711, 8174, 324, -8190, 62, 8187, -449, -8166, 
--834, 8126, -1220, -8069, 1600, 7992, -1980, -7900, 2353, 7787, -2723, -7659, 3085, 7512, -3442, -7350, 3790, 7169, -4131, -6974, 4461, 6761, -4783, -6534, 5093, 6291, -5393, -6036, 5680, 5764, 
---5955, -5482, 6215, 5184, -6463, -4877, 6695, 4557, -6913, -4228, 7114, 3887, -7301, -3539, 7469, 3181, -7622, -2818, 7756, 2446, -7874, -2070, 7972, 1687, -8054, -1302, 8115, 912, -8160, -522, 
--8184, 128, -8191, 265, 8177, -658, -8147, 1049, 8095, -1439, -8027, 1824, 7938, -2208, -7833, 2584, 7708, -2956, -7566, 3320, 7405, -3678, -7229, 4026, 7033, -4366, -6823, 4695, 6596, -5015, 
---6354, 5321, 6096, -5617, -5825, 5898, 5539, -6167, -5241, 6420, 4929, -6660, -4607, 6882, 4272, -7091, -3929, 7280, 3574, -7455, -3213, 7610, 2842, -7749, -2466, 7868, 2083, -7971, -1696, 8052, 
--1303, -8117, -908, 8160, 509, -8186, -111, 8190, -290, -8177, 688, 8142, -1087, -8090, 1481, 8017, -1874, -7926, 2261, 7815, -2644, -7686, 3019, 7537, -3390, -7372, 3750, 7187, -4103, -6987, 
--4445, 6768, -4778, -6534, 5098, 6283, -5408, -6018, 5703, 5737, -5986, -5443, 6253, 5134, -6507, -4815, 6743, 4482, -6965, -4140, 7168, 3785, -7355, -3423, 7523, 3051, -7675, -2673, 7806, 2286, 
---7920, -1896, 8013, 1498, -8088, -1099, 8141, 695, -8177, -291, 8190, -116, -8185, 521, 8158, -926, -8114, 1328, 8047, -1728, -7962, 2123, 7855, -2514, -7731, 2898, 7586, -3276, -7424, 3645, 
--7242, -4006, -7043, 4356, 6825, -4697, -6592, 5025, 6340, -5342, -6075, 5645, 5792, -5935, -5496, 6208, 5185, -6469, -4863, 6711, 4526, -6938, -4180, 7147, 3821, -7339, -3454, 7511, 3077, -7666, 
---2693, 7800, 2301, -7917, -1905, 8011, 1501, -8088, -1096, 8142, 686, -8177, -276, 8190, -137, -8184, 548, 8156, -960, -8108, 1368, 8038, -1774, -7950, 2174, 7839, -2570, -7711, 2959, 7560, 
---3341, -7392, 3714, 7204, -4079, -6998, 4432, 6773, -4776, -6532, 5105, 6273, -5424, -5999, 5727, 5708, -6018, -5404, 6291, 5084, -6550, -4752, 6790, 4406, -7015, -4051, 7220, 3683, -7408, -3307, 
--7575, 2921, -7725, -2529, 7852, 2128, -7962, -1723, 8049, 1312, -8117, -899, 8161, 482, -8187, -65, 8189, -355, -8172, 771, 8132, -1188, -8072, 1600, 7989, -2009, -7887, 2412, 7763, -2811, 
---7620, 3200, 7455, -3583, -7272, 3955, 7068, -4319, -6848, 4669, 6607, -5010, -6350, 5335, 6075, -5648, -5786, 5945, 5479, -6228, -5159, 6492, 4824, -6742, -4478, 6972, 4117, -7185, -3748, 7377, 
--3366, -7552, -2978, 7705, 2579, -7839, -2175, 7950, 1763, -8042, -1348, 8111, 928, -8160, -506, 8185, 81, -8190, 342, 8172, -766, -8133, 1187, 8070, -1607, -7988, 2020, 7882, -2431, -7757, 
--2833, 7609, -3229, -7442, 3615, 7253, -3993, -7046, 4359, 6818, -4715, -6574, 5056, 6309, -5386, -6029, 5700, 5731, -6000, -5419, 6281, 5090, -6548, -4749, 6795, 4393, -7026, -4027, 7235, 3648, 
---7427, -3260, 7597, 2861, -7748, -2457, 7875, 2043, -7983, -1626, 8068, 1201, -8132, -776, 8171, 346, -8190, 83, 8185, -514, -8159, 942, 8109, -1369, -8038, 1791, 7942, -2210, -7827, 2621, 
--7688, -3027, -7529, 3423, 7348, -3812, -7148, 4188, 6926, -4554, -6686, 4906, 6426, -5247, -6150, 5571, 5855, -5881, -5545, 6174, 5217, -6451, -4876, 6708, 4520, -6948, -4153, 7167, 3772, -7368, 
---3382, 7547, 2981, -7706, -2573, 7842, 2156, -7957, -1734, 8048, 1305, -8119, -874, 8164, 439, -8188, -4, 8188, -433, -8166, 867, 8118, -1300, -8050, 1729, 7957, -2154, -7843, 2572, 7705, 
---2984, -7546, 3386, 7364, -3781, -7163, 4163, 6940, -4535, -6698, 4892, 6435, -5238, -6156, 5566, 5857, -5881, -5542, 6177, 5210, -6458, -4865, 6718, 4503, -6961, -4131, 7181, 3744, -7384, -3348, 
--7563, 2940, -7722, -2526, 7857, 2102, -7971, -1674, 8060, 1239, -8128, -802, 8170, 361, -8190, 80, 8185, -523, -8158, 962, 8105, -1401, -8030, 1834, 7930, -2263, -7809, 2684, 7662, -3100, 
---7496, 3505, 7305, -3901, -7095, 4285, 6862, -4657, -6610, 5015, 6337, -5360, -6047, 5687, 5738, -5999, -5413, 6292, 5070, -6569, -4714, 6824, 4342, -7061, -3959, 7276, 3562, -7471, -3156, 7641, 
--2739, -7792, -2315, 7917, 1882, -8021, -1446, 8098, 1003, -8154, -559, 8184, 111, -8191, 336, 8171, -783, -8130, 1227, 8061, -1669, -7971, 2104, 7855, -2535, -7717, 2957, 7554, -3372, -7370, 
--3775, 7162, -4169, -6934, 4549, 6683, -4917, -6414, 5268, 6124, -5606, -5817, 5925, 5490, -6228, -5149, 6510, 4789, -6774, -4417, 7017, 4030, -7240, -3632, 7439, 3221, -7618, -2801, 7771, 2372, 
---7903, -1936, 8009, 1493, -8092, -1047, 8149, 595, -8183, -144, 8190, -310, -8174, 762, 8131, -1213, -8065, 1659, 7972, -2102, -7856, 2536, 7714, -2965, -7551, 3383, 7362, -3793, -7153, 4189, 
--6919, -4575, -6665, 4944, 6390, -5301, -6096, 5639, 5781, -5962, -5450, 6264, 5100, -6549, -4736, 6812, 4355, -7056, -3963, 7276, 3556, -7476, -3140, 7650, 2711, -7802, -2276, 7928, 1832, -8032, 
---1384, 8108, 930, -8161, -474, 8187, 14, -8189, 443, 8163, -902, -8113, 1355, 8036, -1807, -7936, 2251, 7809, -2691, -7659, 3120, 7482, -3541, -7284, 3950, 7061, -4348, -6818, 4730, 6551, 
---5100, -6265, 5451, 5957, -5788, -5631, 6104, 5286, -6403, -4926, 6680, 4548, -6938, -4158, 7171, 3752, -7384, -3336, 7572, 2907, -7737, -2471, 7876, 2024, -7991, -1573, 8079, 1115, -8144, -655, 
--8180, 190, -8191, 273, 8175, -737, -8134, 1198, 8065, -1656, -7972, 2108, 7851, -2555, -7707, 2992, 7536, -3421, -7343, 3838, 7123, -4244, -6883, 4635, 6618, -5013, -6334, 5372, 6027, -5717, 
---5702, 6041, 5356, -6347, -4995, 6631, 4616, -6896, -4223, 7136, 3814, -7355, -3395, 7548, 2963, -7718, -2522, 7862, 2071, -7981, -1616, 8073, 1152, -8140, -687, 8178, 217, -8191, 251, 8176, 
---721, -8136, 1187, 8067, -1651, -7973, 2108, 7851, -2560, -7704, 3002, 7531, -3436, -7334, 3857, 7111, -4267, -6867, 4662, 6597, -5043, -6308, 5405, 5995, -5752, -5665, 6077, 5313, -6385, -4945, 
--6669, 4559, -6934, -4160, 7173, 3744, -7390, -3318, 7581, 2879, -7749, -2432, 7888, 1974, -8004, -1512, 8090, 1042, -8152, -571, 8184, 95, -8190, 379, 8167, -854, -8119, 1324, 8041, -1792, 
---7938, 2252, 7806, -2707, -7650, 3150, 7465, -3586, -7258, 4007, 7024, -4417, -6767, 4810, 6486, -5189, -6185, 5548, 5860, -5891, -5518, 6212, 5154, -6514, -4775, 6791, 4378, -7048, -3967, 7279, 
--3540, -7487, -3104, 7667, 2654, -7824, -2197, 7951, 1731, -8054, -1260, 8126, 783, -8173, -305, 8190, -176, -8181, 655, 8142, -1134, -8076, 1607, 7981, -2076, -7860, 2537, 7710, -2991, -7535, 
--3433, 7332, -3866, -7105, 4283, 6852, -4687, -6577, 5074, 6277, -5445, -5957, 5795, 5615, -6127, -5254, 6436, 4874, -6724, -4478, 6988, 4064, -7229, -3638, 7443, 3197, -7633, -2747, 7794, 2285, 
---7930, -1816, 8037, 1340, -8117, -860, 8167, 375, -8190, 109, 8183, -596, -8149, 1078, 8084, -1559, -7992, 2032, 7870, -2501, -7723, 2959, 7546, -3408, -7344, 3844, 7115, -4268, -6862, 4675, 
--6583, -5068, -6282, 5441, 5957, -5797, -5612, 6131, 5246, -6445, -4862, 6734, 4459, -7001, -4042, 7241, 3609, -7458, -3165, 7646, 2707, -7809, -2241, 7942, 1765, -8048, -1284, 8124, 797, -8173, 
---308, 8190, -183, -8180, 673, 8139, -1162, -8070, 1645, 7971, -2124, -7844, 2594, 7687, -3056, -7505, 3506, 7293, -3946, -7057, 4369, 6793, -4779, -6507, 5169, 6195, -5543, -5862, 5895, 5506, 
---6228, -5132, 6536, 4737, -6823, -4326, 7082, 3898, -7319, -3457, 7526, 3002, -7709, -2537, 7861, 2061, -7987, -1579, 8081, 1090, -8148, -598, 8183, 101, -8190, 393, 8165, -889, -8113, 1380, 
--8028, -1867, -7916, 2346, 7772, -2819, -7602, 3279, 7402, -3730, -7177, 4165, 6923, -4586, -6645, 4989, 6341, -5376, -6015, 5741, 5664, -6086, -5295, 6408, 4904, -6707, -4496, 6980, 4070, -7229, 
---3630, 7450, 3175, -7644, -2709, 7809, 2232, -7946, -1747, 8052, 1254, -8129, -759, 8175, 258, -8191, 242, 8176, -743, -8131, 1240, 8054, -1734, -7949, 2220, 7812, -2700, -7648, 3168, 7452, 
---3626, -7231, 4068, 6980, -4498, -6705, 4908, 6403, -5303, -6078, 5675, 5728, -6028, -5359, 6357, 4967, -6663, -4558, 6943, 4129, -7198, -3687, 7424, 3229, -7624, -2760, 7793, 2278, -7935, -1790, 
--8044, 1292, -8125, -792, 8173, 286, -8191, 219, 8177, -725, -8133, 1227, 8056, -1726, -7950, 2217, 7812, -2701, -7646, 3174, 7448, -3636, -7224, 4083, 6970, -4516, -6691, 4930, 6384, -5327, 
---6055, 5702, 5700, -6057, -5325, 6386, 4927, -6693, -4512, 6973, 4078, -7227, -3629, 7452, 3164, -7650, -2689, 7817, 2202, -7955, -1707, 8060, 1204, -8136, -698, 8179, 187, -8191, 323, 8170, 
---834, -8119, 1340, 8034, -1843, -7920, 2337, 7773, -2824, -7598, 3298, 7390, -3761, -7156, 4208, 6892, -4640, -6602, 5053, 6285, -5447, -5944, 5819, 5578, -6170, -5193, 6494, 4784, -6796, -4359, 
--7068, 3914, -7315, -3455, 7531, 2981, -7719, -2497, 7875, 2001, -8002, -1498, 8096, 988, -8159, -475, 8188, -41, -8186, 556, 8150, -1071, -8084, 1579, 7983, -2084, -7853, 2578, 7689, -3064, 
---7496, 3537, 7272, -3997, -7020, 4440, 6739, -4867, -6432, 5273, 6098, -5659, -5741, 6022, 5358, -6362, -4956, 6675, 4533, -6963, -4092, 7221, 3634, -7453, -3162, 7652, 2675, -7823, -2180, 7960, 
--1673, -8068, -1162, 8141, 644, -8182, -125, 8189, -397, -8165, 915, 8106, -1432, -8016, 1942, 7891, -2445, -7736, 2937, 7548, -3419, -7331, 3885, 7082, -4338, -6807, 4771, 6501, -5187, -6171, 
--5580, 5814, -5953, -5434, 6299, 5031, -6622, -4608, 6915, 4165, -7183, -3706, 7419, 3231, -7627, -2743, 7802, 2242, -7946, -1734, 8056, 1217, -8135, -696, 8179, 170, -8191, 354, 8167, -880, 
---8112, 1400, 8021, -1916, -7899, 2423, 7742, -2922, -7555, 3406, 7335, -3879, -7086, 4335, 6806, -4774, -6500, 5192, 6164, -5590, -5805, 5963, 5419, -6313, -5013, 6636, 4584, -6933, -4138, 7199, 
--3672, -7437, -3192, 7642, 2697, -7818, -2193, 7958, 1677, -8068, -1156, 8142, 628, -8183, -100, 8189, -432, -8162, 960, 8099, -1486, -8003, 2003, 7872, -2515, -7710, 3014, 7514, -3503, -7287, 
--3975, 7028, -4433, -6741, 4870, 6424, -5288, -6081, 5683, 5710, -6055, -5317, 6400, 4899, -6720, -4463, 7010, 4005, -7272, -3532, 7501, 3042, -7701, -2541, 7865, 2027, -7999, -1506, 8096, 977, 
---8161, -445, 8189, -91, -8184, 625, 8142, -1159, -8067, 1685, 7956, -2207, -7812, 2717, 7633, -3218, -7424, 3703, 7180, -4175, -6908, 4626, 6603, -5060, -6272, 5471, 5912, -5860, -5529, 6222, 
--5119, -6559, -4690, 6866, 4237, -7145, -3769, 7392, 3282, -7609, -2782, 7791, 2269, -7941, -1747, 8055, 1215, -8136, -680, 8180, 140, -8190, 398, 8163, -938, -8102, 1471, 8004, -2001, -7873, 
--2519, 7706, -3029, -7507, 3524, 7273, -4006, -7009, 4468, 6713, -4913, -6389, 5335, 6035, -5735, -5656, 6109, 5250, -6458, -4824, 6776, 4374, -7067, -3906, 7325, 3419, -7553, -2919, 7745, 2404, 
---7906, -1880, 8030, 1346, -8120, -808, 8173, 263, -8191, 280, 8172, -825, -8118, 1364, 8026, -1899, -7901, 2424, 7738, -2941, -7543, 3442, 7313, -3931, -7052, 4400, 6758, -4852, -6435, 5280, 
--6081, -5687, -5703, 6067, 5297, -6422, -4869, 6746, 4417, -7042, -3947, 7305, 3457, -7537, -2954, 7734, 2435, -7898, -1908, 8025, 1369, -8118, -826, 8172, 277, -8191, 271, 8172, -820, -8118, 
--1364, 8026, -1903, -7899, 2433, 7735, -2953, -7537, 3459, 7304, -3951, -7039, 4423, 6741, -4878, -6413, 5308, 6055, -5717, -5671, 6098, 5260, -6453, -4826, 6777, 4368, -7073, -3892, 7334, 3396, 
---7564, -2887, 7758, 2362, -7919, -1829, 8041, 1285, -8129, -736, 8178, 183, -8191, 370, 8165, -923, -8103, 1471, 8003, -2013, -7868, 2545, 7694, -3067, -7487, 3574, 7244, -4066, -6970, 4537, 
--6661, -4990, -6323, 5418, 5955, -5823, -5560, 6200, 5138, -6550, -4694, 6868, 4226, -7156, -3741, 7410, 3236, -7631, -2718, 7815, 2185, -7964, -1643, 8075, 1092, -8151, -538, 8186, -21, -8186, 
--578, 8146, -1135, -8069, 1684, 7953, -2228, -7802, 2760, 7613, -3281, -7390, 3785, 7130, -4273, -6839, 4739, 6514, -5186, -6160, 5606, 5775, -6003, -5365, 6369, 4928, -6708, -4470, 7013, 3988, 
---7287, -3489, 7526, 2972, -7730, -2443, 7897, 1900, -8028, -1350, 8120, 791, -8176, -231, 8190, -333, -8168, 894, 8106, -1452, -8007, 2002, 7868, -2545, -7694, 3073, 7482, -3590, -7235, 4087, 
--6953, -4567, -6639, 5024, 6292, -5459, -5916, 5866, 5510, -6247, -5080, 6597, 4624, -6917, -4147, 7203, 3648, -7456, -3134, 7671, 2602, -7852, -2060, 7994, 1506, -8099, -947, 8164, 380, -8191, 
--186, 8177, -754, -8126, 1316, 8034, -1874, -7905, 2421, 7736, -2959, -7531, 3480, 7289, -3988, -7013, 4474, 6701, -4940, -6359, 5381, 5984, -5798, -5581, 6185, 5150, -6545, -4696, 6871, 4216, 
---7165, -3719, 7423, 3200, -7647, -2669, 7832, 2122, -7981, -1566, 8089, 1001, -8160, -432, 8189, -140, -8180, 711, 8130, -1279, -8041, 1840, 7912, -2394, -7745, 2935, 7539, -3463, -7298, 3973, 
--7019, -4465, -6707, 4934, 6361, -5380, -5985, 5799, 5577, -6191, -5144, 6550, 4684, -6880, -4202, 7174, 3698, -7434, -3177, 7656, 2638, -7843, -2088, 7988, 1526, -8097, -958, 8163, 383, -8191, 
--192, 8176, -769, -8123, 1340, 8028, -1906, -7895, 2461, 7720, -3006, -7509, 3534, 7259, -4047, -6975, 4538, 6654, -5009, -6301, 5453, 5915, -5871, -5502, 6259, 5058, -6617, -4592, 6941, 4100, 
---7232, -3590, 7485, 3059, -7702, -2515, 7879, 1956, -8019, -1389, 8116, 814, -8175, -235, 8190, -346, -8167, 924, 8100, -1500, -7995, 2066, 7847, -2624, -7662, 3167, 7436, -3697, -7174, 4205, 
--6874, -4695, -6542, 5159, 6174, -5599, -5776, 6009, 5348, -6391, -4894, 6738, 4413, -7054, -3912, 7331, 3388, -7574, -2849, 7776, 2294, -7940, -1728, 8063, 1152, -8146, -572, 8186, -14, -8186, 
--598, 8142, -1180, -8059, 1755, 7932, -2324, -7767, 2878, 7560, -3420, -7316, 3943, 7033, -4447, -6716, 4927, 6362, -5384, -5977, 5811, 5559, -6211, -5115, 6577, 4642, -6911, -4148, 7207, 3629, 
---7469, -3094, 7690, 2541, -7874, -1976, 8015, 1399, -8116, -816, 8174, 227, -8191, 361, 8164, -949, -8097, 1531, 7986, -2108, -7835, 2671, 7641, -3223, -7410, 3756, 7138, -4272, -6831, 4763, 
--6487, -5232, -6110, 5672, 5699, -6085, -5261, 6464, 4793, -6811, -4302, 7121, 3786, -7396, -3252, 7630, 2699, -7826, -2134, 7980, 1555, -8094, -970, 8163, 378, -8191, 215, 8174, -809, -8117, 
--1396, 8015, -1978, -7872, 2549, 7686, -3107, -7462, 3648, 7196, -4172, -6894, 4672, 6553, -5149, -6180, 5597, 5772, -6018, -5335, 6405, 4868, -6760, -4377, 7078, 3861, -7360, -3326, 7601, 2771, 
---7804, -2203, 7964, 1621, -8083, -1033, 8157, 437, -8190, 160, 8178, -758, -8123, 1350, 8024, -1937, -7883, 2512, 7698, -3076, -7475, 3622, 7209, -4150, -6906, 4654, 6564, -5136, -6189, 5588, 
--5779, -6012, -5340, 6403, 4870, -6760, -4375, 7080, 3855, -7364, -3316, 7606, 2757, -7810, -2184, 7969, 1598, -8087, -1005, 8160, 405, -8191, 196, 8175, -798, -8118, 1394, 8014, -1985, -7869, 
--2563, 7679, -3129, -7450, 3677, 7178, -4207, -6869, 4712, 6521, -5194, -6139, 5645, 5722, -6068, -5275, 6456, 4798, -6812, -4296, 7128, 3768, -7407, -3222, 7644, 2656, -7841, -2078, 7994, 1486, 
---8105, -887, 8170, 282, -8191, 323, 8166, -929, -8099, 1528, 7985, -2120, -7828, 2699, 7627, -3266, -7386, 3813, 7102, -4341, -6781, 4843, 6421, -5320, -6027, 5767, 5598, -6184, -5139, 6565, 
--4650, -6911, -4138, 7218, 3600, -7487, -3044, 7712, 2469, -7897, -1882, 8036, 1283, -8132, -678, 8182, 68, -8188, 541, 8147, -1150, -8062, 1750, 7930, -2343, -7757, 2921, 7538, -3484, -7279, 
--4027, 6977, -4549, -6638, 5044, 6260, -5513, -5849, 5949, 5403, -6354, -4929, 6722, 4425, -7054, -3898, 7345, 3347, -7597, -2779, 7804, 2193, -7969, -1597, 8088, 989, -8163, -378, 8190, -237, 
---8173, 850, 8109, -1460, -8000, 2059, 7844, -2650, -7646, 3223, 7403, -3781, -7120, 4315, 6794, -4827, -6432, 5310, 6032, -5765, -5599, 6185, 5132, -6573, -4638, 6921, 4115, -7232, -3571, 7501, 
--3005, -7728, -2423, 7910, 1825, -8049, -1219, 8140, 603, -8186, 14, 8184, -633, -8137, 1247, 8042, -1856, -7903, 2452, 7716, -3037, -7488, 3603, 7214, -4150, -6901, 4671, 6546, -5168, -6156, 
--5633, 5728, -6068, -5269, 6466, 4778, -6830, -4261, 7152, 3717, -7435, -3154, 7673, 2570, -7870, -1974, 8018, 1364, -8123, -748, 8179, 125, -8189, 497, 8151, -1118, -8067, 1730, 7934, -2335, 
---7757, 2925, 7533, -3499, -7268, 4052, 6958, -4583, -6610, 5086, 6221, -5562, -5798, 6003, 5339, -6411, -4851, 6780, 4332, -7112, -3790, 7400, 3224, -7648, -2641, 7849, 2040, -8006, -1429, 8114, 
--807, -8177, -183, 8189, -445, -8156, 1068, 8074, -1688, -7945, 2295, 7769, -2891, -7548, 3469, 7281, -4028, -6973, 4562, 6622, -5071, -6234, 5548, 5807, -5995, -5348, 6405, 4855, -6779, -4335, 
--7111, 3788, -7403, -3220, 7650, 2630, -7853, -2027, 8008, 1410, -8117, -786, 8177, 156, -8190, 474, 8152, -1103, -8068, 1724, 7935, -2337, -7755, 2934, 7528, -3515, -7258, 4074, 6942, -4611, 
---6588, 5119, 6191, -5598, -5760, 6042, 5292, -6452, -4794, 6822, 4266, -7152, -3714, 7439, 3137, -7682, -2544, 7878, 1933, -8029, -1312, 8130, 681, -8183, -48, 8186, -587, -8142, 1218, 8046, 
---1843, -7904, 2455, 7713, -3055, -7477, 3634, 7193, -4194, -6869, 4726, 6501, -5232, -6095, 5705, 5650, -6145, -5174, 6547, 4663, -6910, -4127, 7231, 3563, -7509, -2979, 7740, 2375, -7926, -1759, 
--8062, 1130, -8151, -495, 8189, -144, -8178, 781, 8116, -1416, -8007, 2040, 7847, -2653, -7641, 3249, 7386, -3827, -7088, 4380, 6744, -4908, -6362, 5405, 5938, -5870, -5480, 6298, 4986, -6689, 
---4463, 7037, 3911, -7345, -3337, 7605, 2740, -7821, -2128, 7987, 1501, -8105, -866, 8172, 224, -8191, 418, 8157, -1059, -8075, 1692, 7941, -2317, -7760, 2925, 7529, -3518, -7254, 4087, 6931, 
---4634, -6568, 5149, 6162, -5635, -5719, 6084, 5239, -6498, -4729, 6869, 4186, -7200, -3620, 7484, 3029, -7724, -2421, 7914, 1796, -8057, -1161, 8147, 517, -8189, 128, 8178, -775, -8118, 1415, 
--8005, -2049, -7844, 2668, 7632, -3272, -7375, 3854, 7069, -4414, -6720, 4945, 6328, -5447, -5898, 5913, 5428, -6344, -4927, 6733, 4392, -7083, -3832, 7385, 3245, -7644, -2640, 7852, 2016, -8013, 
---1381, 8122, 735, -8181, -87, 8187, -565, -8143, 1211, 8046, -1851, -7900, 2478, 7702, -3092, -7457, 3684, 7163, -4255, -6825, 4797, 6442, -5311, -6020, 5790, 5558, -6234, -5062, 6636, 4532, 
---6998, -3975, 7314, 3391, -7586, -2787, 7807, 2162, -7981, -1526, 8102, 878, -8173, -227, 8190, -429, -8157, 1080, 8069, -1726, -7932, 2359, 7743, -2980, -7505, 3579, 7218, -4158, -6886, 4708, 
--6508, -5231, -6090, 5718, 5631, -6170, -5137, 6581, 4608, -6951, -4052, 7275, 3467, -7554, -2862, 7783, 2236, -7964, -1598, 8091, 947, -8168, -291, 8190, -368, -8162, 1023, 8079, -1674, -7945, 
--2312, 7758, -2937, -7523, 3542, 7236, -4125, -6905, 4680, 6527, -5207, -6109, 5699, 5648, -6155, -5153, 6569, 4622, -6943, -4063, 7270, 3475, -7552, -2867, 7782, 2238, -7964, -1595, 8092, 941, 
---8169, -281, 8190, -382, -8161, 1041, 8075, -1695, -7939, 2336, 7749, -2964, -7510, 3571, 7220, -4157, -6884, 4714, 6501, -5242, -6078, 5733, 5612, -6189, -5111, 6603, 4574, -6975, -4009, 7299, 
--3416, -7578, -2802, 7804, 2167, -7981, -1520, 8103, 860, -8174, -197, 8189, -470, -8152, 1132, 8059, -1789, -7914, 2432, 7715, -3061, -7467, 3668, 7167, -4253, -6822, 4808, 6429, -5333, -5996, 
--5821, 5520, -6272, -5009, 6679, 4463, -7045, -3889, 7361, 3288, -7631, -2665, 7847, 2023, -8014, -1370, 8124, 705, -8183, -37, 8185, -634, -8134, 1298, 8027, -1956, -7868, 2599, 7654, -3227, 
---7391, 3831, 7076, -4412, -6716, 4961, 6308, -5479, -5860, 5958, 5370, -6400, -4846, 6797, 4288, -7149, -3702, 7452, 3089, -7707, -2457, 7908, 1806, -8057, -1145, 8150, 474, -8190, 198, 8173, 
---871, -8102, 1537, 7975, -2194, -7795, 2835, 7561, -3459, -7277, 4057, 6942, -4630, -6561, 5170, 6134, -5676, -5667, 6143, 5160, -6569, -4619, 6949, 4044, -7284, -3444, 7567, 2818, -7801, -2175, 
--7980, 1514, -8106, -845, 8175, 169, -8190, 508, 8147, -1182, -8050, 1847, 7896, -2502, -7690, 3138, 7429, -3754, -7119, 4343, 6758, -4904, -6353, 5429, 5902, -5920, -5412, 6367, 4883, -6773, 
---4322, 7131, 3729, -7442, -3112, 7699, 2472, -7905, -1816, 8055, 1146, -8151, -470, 8189, -212, -8173, 891, 8098, -1565, -7969, 2227, 7782, -2876, -7544, 3503, 7251, -4108, -6910, 4683, 6519, 
---5227, -6084, 5733, 5605, -6201, -5089, 6625, 4535, -7004, -3952, 7333, 3339, -7613, -2704, 7837, 2049, -8010, -1381, 8124, 701, -8184, -18, 8184, -667, -8129, 1346, 8016, -2018, -7848, 2673, 
--7623, -3312, -7347, 3927, 7017, -4515, -6640, 5070, 6214, -5592, -5746, 6073, 5236, -6513, -4691, 6905, 4111, -7251, -3503, 7544, 2869, -7786, -2217, 7971, 1546, -8102, -867, 8174, 179, -8190, 
--509, 8146, -1195, -8047, 1870, 7888, -2535, -7676, 3180, 7407, -3804, -7088, 4400, 6717, -4967, -6299, 5496, 5835, -5989, -5332, 6437, 4788, -6842, -4212, 7196, 3604, -7501, -2972, 7751, 2317, 
---7948, -1647, 8086, 963, -8168, -274, 8190, -419, -8156, 1107, 8061, -1790, -7911, 2458, 7702, -3110, -7440, 3739, 7122, -4343, -6756, 4914, 6339, -5452, -5878, 5948, 5373, -6405, -4831, 6813, 
--4253, -7175, -3645, 7483, 3010, -7739, -2354, 7938, 1679, -8081, -994, 8165, 300, -8191, 395, 8157, -1089, -8065, 1773, 7913, -2447, -7706, 3101, 7442, -3735, -7125, 4341, 6754, -4917, -6337, 
--5455, 5872, -5956, -5365, 6412, 4818, -6824, -4238, 7184, 3624, -7494, -2986, 7747, 2324, -7947, -1648, 8086, 957, -8169, -260, 8190, -440, -8153, 1135, 8055, -1825, -7901, 2499, 7686, -3157, 
---7417, 3790, 7092, -4398, -6717, 4971, 6290, -5511, -5820, 6008, 5304, -6463, -4752, 6869, 4163, -7227, -3544, 7529, 2898, -7779, -2232, 7969, 1548, -8103, -854, 8175, 151, -8189, 551, 8141, 
---1251, -8034, 1939, 7867, -2616, -7643, 3272, 7361, -3906, -7026, 4509, 6637, -5081, -6201, 5613, 5718, -6106, -5193, 6552, 4628, -6951, -4031, 7297, 3401, -7591, -2748, 7827, 2072, -8007, -1383, 
--8125, 682, -8185, 23, 8182, -730, -8120, 1430, 7995, -2121, -7813, 2795, 7571, -3450, -7274, 4077, 6921, -4676, -6518, 5238, 6064, -5764, -5566, 6244, 5025, -6680, -4448, 7064, 3836, -7397, 
---3196, 7673, 2531, -7893, -1848, 8052, 1149, -8153, -444, 8190, -267, -8168, 974, 8082, -1677, -7938, 2364, 7732, -3036, -7469, 3684, 7148, -4306, -6775, 4893, 6349, -5446, -5877, 5955, 5358, 
---6422, -4801, 6839, 4205, -7206, -3579, 7516, 2924, -7772, -2249, 7966, 1554, -8103, -850, 8176, 136, -8189, 576, 8137, -1286, -8026, 1985, 7852, -2671, -7620, 3335, 7328, -3975, -6982, 4584, 
--6581, -5159, -6132, 5694, 5633, -6187, -5094, 6631, 4513, -7026, -3900, 7366, 3255, -7652, -2587, 7877, 1896, -8044, -1194, 8148, 479, -8191, 237, 8169, -953, -8086, 1661, 7940, -2358, -7734, 
--3034, 7467, -3690, -7145, 4316, 6765, -4910, -6335, 5465, 5855, -5980, -5331, 6447, 4763, -6866, -4161, 7231, 3525, -7542, -2863, 7792, 2177, -7985, -1476, 8114, 761, -8182, -43, 8184, -679, 
---8126, 1393, 8002, -2099, -7818, 2786, 7572, -3454, -7268, 4094, 6907, -4704, -6493, 5275, 6027, -5808, -5515, 6293, 4959, -6732, -4366, 7116, 3737, -7447, -3080, 7718, 2397, -7931, -1698, 8080, 
--983, -8168, -262, 8190, -464, -8150, 1183, 8044, -1896, -7877, 2592, 7647, -3270, -7358, 3921, 7010, -4543, -6609, 5127, 6154, -5674, -5652, 6173, 5103, -6627, -4517, 7027, 3892, -7373, -3239, 
--7659, 2559, -7887, -1859, 8051, 1143, -8154, -420, 8190, -309, -8164, 1033, 8071, -1752, -7916, 2454, 7697, -3140, -7419, 3799, 7080, -4430, -6686, 5024, 6238, -5581, -5742, 6091, 5199, -6555, 
---4616, 6966, 3994, -7323, -3342, 7619, 2662, -7858, -1962, 8032, 1244, -8144, -518, 8189, -214, -8171, 942, 8086, -1666, -7938, 2374, 7725, -3065, -7452, 3730, 7118, -4368, -6728, 4968, 6283, 
---5531, -5789, 6048, 5246, -6519, -4664, 6935, 4042, -7298, -3389, 7601, 2707, -7845, -2005, 8023, 1285, -8139, -556, 8188, -179, -8173, 911, 8090, -1638, -7944, 2350, 7732, -3046, -7460, 3715, 
--7125, -4356, -6735, 4960, 6288, -5526, -5792, 6046, 5248, -6519, -4663, 6937, 4037, -7302, -3381, 7605, 2696, -7849, -1990, 8027, 1266, -8142, -534, 8189, -205, -8171, 940, 8086, -1670, -7936, 
--2385, 7720, -3083, -7443, 3753, 7103, -4395, -6707, 5000, 6255, -5565, -5753, 6084, 5203, -6555, -4611, 6971, 3980, -7332, -3319, 7631, 2627, -7869, -1917, 8042, 1188, -8150, -451, 8190, -291, 
---8165, 1029, 8071, -1761, -7912, 2477, 7686, -3175, -7400, 3845, 7050, -4485, -6644, 5087, 6182, -5648, -5671, 6162, 5110, -6627, -4510, 7035, 3870, -7388, -3200, 7677, 2501, -7906, -1784, 8067, 
--1050, -8163, -308, 8190, -438, -8151, 1178, 8043, -1911, -7870, 2626, 7630, -3322, -7329, 3988, 6964, -4624, -6544, 5219, 6068, -5773, -5542, 6277, 4969, -6732, -4356, 7128, 3705, -7467, -3024, 
--7742, 2317, -7954, -1592, 8099, 851, -8178, -105, 8186, -644, -8128, 1386, 8001, -2118, -7808, 2831, 7548, -3523, -7227, 4183, 6843, -4810, -6404, 5395, 5909, -5937, -5366, 6428, 4776, -6866, 
---4148, 7245, 3483, -7566, -2791, 7820, 2073, -8012, -1339, 8133, 592, -8189, 159, 8173, -910, -8091, 1652, 7938, -2382, -7720, 3090, 7435, -3774, -7089, 4425, 6682, -5040, -6219, 5611, 5702, 
---6136, -5139, 6608, 4530, -7026, -3884, 7383, 3203, -7679, -2497, 7907, 1768, -8071, -1025, 8165, 271, -8191, 483, 8145, -1235, -8032, 1975, 7849, -2700, -7601, 3400, 7286, -4074, -6911, 4711, 
--6475, -5310, -5986, 5862, 5443, -6366, -4856, 6814, 4225, -7205, -3560, 7533, 2862, -7799, -2142, 7996, 1401, -8127, -649, 8186, -110, -8177, 866, 8096, -1617, -7947, 2352, 7728, -3069, -7445, 
--3758, 7095, -4417, -6686, 5036, 6218, -5614, -5698, 6142, 5127, -6619, -4514, 7037, 3859, -7397, -3173, 7690, 2458, -7920, -1723, 8079, 971, -8170, -212, 8189, -551, -8139, 1307, 8016, -2054, 
---7826, 2781, 7566, -3486, -7242, 4160, 6854, -4799, -6408, 5395, 5904, -5947, -5351, 6444, 4749, -6888, -4108, 7270, 3428, -7591, -2721, 7844, 1988, -8031, -1239, 8145, 478, -8191, 286, 8163, 
---1050, -8066, 1803, 7897, -2542, -7660, 3257, 7354, -3946, -6986, 4598, 6555, -5213, -6068, 5780, 5526, -6298, -4938, 6759, 4304, -7163, -3634, 7503, 2930, -7778, -2202, 7984, 1452, -8121, -692, 
--8185, -77, -8179, 843, 8098, -1604, -7949, 2350, 7727, -3076, -7439, 3774, 7084, -4440, -6668, 5066, 6191, -5649, -5661, 6180, 5079, -6658, -4453, 7076, 3787, -7434, -3088, 7723, 2360, -7946, 
---1613, 8097, 850, -8178, -80, 8185, -692, -8121, 1456, 7982, -2210, -7775, 2942, 7497, -3650, -7153, 4324, 6744, -4961, -6277, 5553, 5752, -6097, -5177, 6584, 4554, -7016, -3893, 7382, 3194, 
---7685, -2469, 7918, 1719, -8081, -956, 8171, 182, -8189, 592, 8132, -1362, -8004, 2119, 7802, -2859, -7533, 3571, 7193, -4254, -6791, 4896, 6326, -5497, -5806, 6046, 5232, -6543, -4612, 6980, 
--3949, -7356, -3252, 7663, 2524, -7904, -1774, 8071, 1007, -8168, -232, 8189, -547, -8138, 1319, 8012, -2082, -7815, 2824, 7545, -3543, -7209, 4227, 6806, -4876, -6343, 5479, 5820, -6034, -5247, 
--6532, 4624, -6974, -3960, 7350, 3259, -7662, -2530, 7902, 1775, -8072, -1007, 8167, 227, -8190, 554, 8136, -1331, -8010, 2095, 7809, -2841, -7539, 3560, 7198, -4249, -6793, 4897, 6324, -5502, 
---5799, 6056, 5219, -6556, -4593, 6994, 3923, -7370, -3218, 7677, 2483, -7916, -1726, 8080, 951, -8172, -169, 8187, -616, -8129, 1394, 7995, -2161, -7789, 2907, 7509, -3628, -7162, 4314, 6747, 
---4963, -6272, 5563, 5737, -6115, -5151, 6609, 4515, -7043, -3839, 7411, 3126, -7713, -2386, 7941, 1622, -8098, -844, 8178, 57, -8185, 730, 8113, -1511, -7969, 2277, 7749, -3024, -7458, 3742, 
--7097, -4426, -6672, 5068, 6182, -5665, -5637, 6207, 5038, -6694, -4393, 7117, 3706, -7475, -2986, 7762, 2236, -7979, -1467, 8120, 682, -8186, 108, 8175, -899, -8089, 1679, 7926, -2446, -7691, 
--3189, 7381, -3903, -7005, 4580, 6561, -5216, -6057, 5801, 5495, -6333, -4883, 6805, 4223, -7215, -3525, 7555, 2792, -7827, -2035, 8023, 1256, -8146, -467, 8190, -328, -8159, 1118, 8050, -1900, 
---7867, 2663, 7607, -3402, -7278, 4108, 6878, -4777, -6415, 5399, 5890, -5972, -5310, 6487, 4679, -6943, -4005, 7331, 3291, -7652, -2547, 7899, 1778, -8073, -993, 8169, 197, -8189, 599, 8130, 
---1392, -7995, 2170, 7783, -2929, -7498, 3659, 7140, -4356, -6717, 5010, 6227, -5618, -5680, 6172, 5077, -6668, -4427, 7099, 3733, -7465, -3005, 7757, 2247, -7978, -1468, 8120, 674, -8187, 125, 
--8174, -925, -8084, 1715, 7915, -2490, -7673, 3240, 7355, -3961, -6968, 4642, 6513, -5280, -5997, 5866, 5421, -6399, -4795, 6867, 4121, -7272, -3410, 7605, 2663, -7868, -1892, 8052, 1102, -8161, 
---302
 
(2459, 563, -2410, -372, 2370, 182, -2321, -1, 2264, 
-184, -2224, 372, 2173, -544, -2126, 724, 2083, -892, 
-2035, 1045, 2001, -1201, -1959, 1355, 1941, -1491, -1900, 
1611, 1887, -1745, -1873, 1847, 1855, -1958, -1851, 2052, 
1836, -2133, -1849, 2217, 1848, -2280, -1851, 2338, 1864, 
-2381, -1892, 2404, 1911, -2432, -1932, 2457, 1953, -2459, 
-1990, 2456, 2014, -2444, -2052, 2424, 2078, -2401, -2112, 
2361, 2157, -2317, -2184, 2262, 2227, -2195, -2251, 2127, 
2299, -2062, -2332, 1979, 2361, -1894, -2375, 1813, 2412, 
-1731, -2432, 1626, 2445, -1546, -2471, 1436, 2483, -1342, 
-2493, 1251, 2499, -1145, -2509, 1066, 2517, -963, -2519, 
873, 2502, -787, -2507, 705, 2504, -618, -2489, 546, 
2479, -474, -2470, 407, 2460, -364, -2447, 314, 2424, 
-269, -2417, 235, 2392, -214, -2382, 195, 2383, -189, 
-2369, 187, 2363, -206, -2358, 233, 2353, -256, -2360, 
303, 2362, -352, -2371, 415, 2378, -482, -2395, 559, 
2422, -641, -2446, 751, 2468, -846, -2502, 969, 2542, 
-1087, -2572, 1210, 2608, -1333, -2658, 1469, 2701, -1609, 
-2761, 1760, 2814, -1908, -2863, 2057, 2906, -2210, -2960, 
2345, 3020, -2500, -3072, 2638, 3126, -2778, -3176, 2920, 
3216, -3064, -3262, 3176, 3304, -3308, -3341, 3417, 3358, 
-3510, -3393, 3601, 3400, -3692, -3418, 3763, 3404, -3819, 
-3407, 3869, 3389, -3899, -3373, 3914, 3333, -3908, -3288, 
3909, 3248, -3874, -3180, 3838, 3112, -3778, -3033, 3696, 
2941, -3614, -2835, 3507, 2728, -3371, -2608, 3247, 2479, 
-3084, -2353, 2932, 2215, -2751, -2068, 2556, 1906, -2364, 
-1750, 2148, 1582, -1933, -1414, 1693, 1245, -1462, -1070, 
1220, 900, -961, -728, 713, 551, -459, -377, 212, 
220, 50, -54, -297, -117, 543, 264, -777, -417, 
1016, 550, -1240, -683, 1464, 819, -1675, -934, 1870, 
1044, -2037, -1137, 2216, 1209, -2364, -1298, 2497, 1349, 
-2611, -1394, 2707, 1438, -2785, -1472, 2845, 1481, -2879, 
-1474, 2885, 1474, -2884, -1449, 2850, 1417, -2806, -1379, 
2724, 1320, -2644, -1262, 2529, 1193, -2386, -1121, 2244, 
1029, -2068, -940, 1887, 838, -1683, -735, 1450, 630, 
-1218, -524, 972, 410, -708, -304, 449, 190, -167, 
-84, -120, -31, 399, 122, -698, -226, 992, 322, 
-1267, -406, 1555, 498, -1843, -577, 2124, 647, -2391, 
-705, 2646, 761, -2898, -801, 3134, 836, -3345, -861, 
3555, 884, -3737, -892, 3888, 892, -4036, -884, 4161, 
854, -4249, -825, 4331, 793, -4380, -743, 4395, 697, 
-4390, -633, 4375, 568, -4322, -498, 4240, 430, -4133, 
-352, 3992, 265, -3841, -188, 3664, 90, -3443, -7, 
3230, -79, -2965, 165, 2705, -237, -2417, 316, 2103, 
-405, -1785, 468, 1435, -535, -1094, 602, 721, -661, 
-356, 708, -35, -750, 420, 791, -802, -819, 1191, 
853, -1596, -866, 1976, 875, -2371, -875, 2744, 855, 
-3111, -839, 3481, 828, -3831, -804, 4175, 763, -4484, 
-721, 4796, 684, -5085, -627, 5365, 570, -5618, -522, 
5851, 459, -6055, -399, 6237, 341, -6411, -281, 6557, 
221, -6672, -161, 6768, 107, -6840, -63, 6892, 14, 
-6912, 29, 6914, -65, -6904, 107, 6867, -126, -6809, 
148, 6727, -152, -6633, 166, 6522, -166, -6385, 142, 
6237, -129, -6089, 97, 5925, -64, -5753, 18, 5561, 
20, -5365, -77, 5178, 145, -4974, -227, 4773, 303, 
-4555, -375, 4364, 462, -4161, -548, 3961, 636, -3775, 
-738, 3591, 830, -3412, -911, 3259, 1009, -3094, -1093, 
2949, 1179, -2817, -1266, 2703, 1328, -2597, -1400, 2498, 
1455, -2419, -1521, 2355, 1563, -2305, -1590, 2261, 1620, 
-2244, -1634, 2237, 1621, -2236, -1616, 2267, 1585, -2293, 
-1558, 2346, 1504, -2391, -1431, 2465, 1351, -2536, -1268, 
2619, 1162, -2713, -1047, 2810, 922, -2906, -783, 3016, 
624, -3112, -462, 3222, 302, -3339, -110, 3438, -68, 
-3536, 266, 3639, -460, -3739, 663, 3833, -867, -3910, 
1066, 3986, -1281, -4041, 1483, 4105, -1687, -4151, 1894, 
4180, -2077, -4201, 2268, 4204, -2452, -4197, 2619, 4180, 
-2796, -4139, 2943, 4091, -3098, -4022, 3230, 3959, -3339, 
-3864, 3451, 3753, -3543, -3636, 3616, 3522, -3687, -3377, 
3733, 3229, -3772, -3061, 3801, 2894, -3793, -2723, 3793, 
2531, -3783, -2344, 3753, 2146, -3710, -1932, 3645, 1732, 
-3587, -1534, 3504, 1323, -3421, -1126, 3334, 915, -3246, 
-720, 3151, 518, -3044, -335, 2947, 152, -2836, 29, 
2732, -180, -2621, 348, 2536, -485, -2441, 624, 2352, 
-750, -2269, 862, 2200, -954, -2135, 1040, 2077, -1096, 
-2037, 1159, 2011, -1191, -1984, 1231, 1979, -1237, -2003, 
1232, 2014, -1209, -2059, 1178, 2102, -1131, -2177, 1081, 
2250, -1013, -2340, 933, 2439, -846, -2559, 753, 2691, 
-635, -2824, 525, 2969, -395, -3122, 275, 3279, -144, 
-3442, 2, 3601, 136, -3779, -264, 3937, 413, -4109, 
-547, 4276, 690, -4442, -810, 4595, 946, -4743, -1063, 
4877, 1186, -5008, -1285, 5127, 1380, -5224, -1475, 5296, 
1552, -5372, -1618, 5424, 1679, -5453, -1728, 5446, 1748, 
-5445, -1775, 5405, 1779, -5353, -1765, 5260, 1748, -5158, 
-1719, 5039, 1668, -4886, -1599, 4708, 1526, -4501, -1444, 
4291, 1346, -4048, -1229, 3774, 1102, -3505, -969, 3200, 
818, -2886, -666, 2536, 490, -2200, -314, 1833, 139, 
-1464, 58, 1085, -243, -680, 451, 298, -650, 110, 
859, -508, -1062, 895, 1274, -1297, -1478, 1684, 1698, 
-2073, -1896, 2443, 2105, -2800, -2313, 3154, 2511, -3479, 
-2690, 3807, 2890, -4096, -3063, 4375, 3245, -4646, -3411, 
4880, 3569, -5096, -3714, 5283, 3852, -5449, -3988, 5583, 
4118, -5695, -4221, 5773, 4332, -5844, -4413, 5872, 4501, 
-5880, -4562, 5865, 4631, -5811, -4675, 5750, 4716, -5660, 
-4734, 5540, 4748, -5400, -4750, 5242, 4734, -5075, -4728, 
4881, 4699, -4670, -4663, 4442, 4606, -4213, -4550, 3955, 
4485, -3711, -4403, 3447, 4319, -3169, -4222, 2896, 4119, 
-2626, -4007, 2353, 3891, -2074, -3760, 1809, 3617, -1535, 
-3478, 1282, 3325, -1032, -3181, 796, 3007, -567, -2849, 
342, 2675, -125, -2482, -62, 2303, 249, -2108, -409, 
1920, 572, -1718, -698, 1520, 816, -1297, -927, 1095, 
1025, -876, -1088, 647, 1148, -430, -1191, 214, 1223, 
14, -1249, -252, 1246, 478, -1236, -710, 1230, 937, 
-1202, -1176, 1161, 1414, -1105, -1643, 1067, 1864, -1001, 
-2095, 942, 2321, -879, -2548, 807, 2766, -749, -2982, 
675, 3179, -602, -3394, 544, 3589, -473, -3784, 427, 
3967, -361, -4139, 327, 4300, -278, -4448, 244, 4608, 
-215, -4744, 197, 4863, -194, -4969, 200, 5075, -201, 
-5161, 221, 5216, -236, -5278, 282, 5322, -315, -5355, 
379, 5368, -427, -5358, 500, 5349, -577, -5317, 659, 
5260, -735, -5211, 823, 5118, -933, -5036, 1023, 4927, 
-1126, -4808, 1236, 4669, -1348, -4512, 1444, 4363, -1564, 
-4189, 1656, 4001, -1775, -3808, 1876, 3603, -1979, -3378, 
2066, 3166, -2163, -2936, 2247, 2703, -2335, -2455, 2410, 
2226, -2490, -1985, 2562, 1729, -2628, -1484, 2684, 1253, 
-2727, -1006, 2762, 771, -2813, -538, 2840, 308, -2870, 
-103, 2885, -107, -2904, 314, 2903, -506, -2913, 683, 
2911, -859, -2916, 1015, 2915, -1154, -2898, 1286, 2883, 
-1403, -2875, 1499, 2874, -1592, -2860, 1662, 2833, -1720, 
-2823, 1758, 2814, -1787, -2798, 1807, 2799, -1806, -2794, 
1790, 2788, -1763, -2788, 1721, 2783, -1671, -2787, 1615, 
2792, -1550, -2800, 1469, 2801, -1379, -2819, 1283, 2829, 
-1183, -2839, 1083, 2850, -977, -2867, 861, 2888, -743, 
-2907, 629, 2932, -522, -2937, 421, 2959, -313, -2970, 
208, 2968, -123, -2971, 39, 2974, 38, -2979, -120, 
2965, 167, -2937, -222, 2926, 263, -2888, -297, 2844, 
306, -2795, -307, 2742, 295, -2671, -276, 2590, 236, 
-2505, -201, 2405, 125, -2290, -55, 2167, -26, -2031, 
110, 1892, -225, -1747, 341, 1577, -463, -1421, 600, 
1237, -741, -1047, 884, 861, -1040, -655, 1195, 446, 
-1346, -242, 1508, 27, -1663, 187, 1829, -407, -1982, 
631, 2130, -847, -2273, 1057, 2411, -1284, -2546, 1481, 
2680, -1692, -2784, 1884, 2884, -2073, -2979, 2243, 3059, 
-2417, -3132, 2567, 3174, -2719, -3216, 2837, 3234, -2946, 
-3233, 3058, 3220, -3128, -3186, 3201, 3142, -3241, -3074, 
3269, 2996, -3283, -2916, 3275, 2790, -3248, -2678, 3191, 
2540, -3127, -2377, 3043, 2225, -2937, -2047, 2819, 1860, 
-2668, -1667, 2510, 1464, -2340, -1253, 2149, 1036, -1942, 
-820, 1718, 592, -1495, -374, 1251, 152, -992, 64, 
733, -273, -462, 489, 186, -692, 84, 881, -373, 
-1068, 653, 1239, -934, -1404, 1218, 1554, -1502, -1688, 
1766, 1804, -2050, -1906, 2302, 1989, -2571, -2055, 2814, 
2113, -3037, -2140, 3261, 2154, -3471, -2150, 3681, 2112, 
-3853, -2069, 4018, 2018, -4175, -1927, 4299, 1833, -4425, 
-1720, 4520, 1596, -4607, -1443, 4661, 1291, -4716, -1126, 
4734, 943, -4745, -745, 4739, 532, -4707, -326, 4653, 
115, -4600, 108, 4527, -326, -4431, 557, 4313, -781, 
-4194, 1001, 4069, -1224, -3911, 1439, 3757, -1655, -3587, 
1848, 3402, -2041, -3216, 2224, 3007, -2398, -2807, 2554, 
2604, -2690, -2392, 2833, 2169, -2943, -1942, 3046, 1718, 
-3123, -1491, 3178, 1258, -3227, -1038, 3258, 817, -3273, 
-590, 3262, 374, -3235, -153, 3186, -64, -3122, 265, 
3051, -466, -2964, 675, 2849, -860, -2733, 1050, 2598, 
-1226, -2443, 1384, 2274, -1562, -2106, 1715, 1930, -1859, 
-1743, 1987, 1548, -2129, -1348, 2249, 1138, -2350, -947, 
2451, 731, -2550, -536, 2638, 331, -2710, -124, 2775, 
-79, -2828, 269, 2875, -460, -2914, 635, 2939, -806, 
-2949, 968, 2957, -1115, -2963, 1258, 2951, -1390, -2920, 
1505, 2896, -1608, -2856, 1699, 2798, -1789, -2734, 1848, 
2669, -1904, -2582, 1947, 2489, -1978, -2386, 1993, 2267, 
-1992, -2143, 1998, 2013, -1979, -1875, 1949, 1722, -1915, 
-1556, 1882, 1383, -1833, -1202, 1762, 1019, -1702, -819, 
1638, 617, -1571, -398, 1493, 167, -1423, 49, 1333, 
-292, -1272, 529, 1188, -780, -1111, 1017, 1051, -1275, 
-985, 1535, 909, -1792, -853, 2045, 802, -2301, -753, 
2565, 714, -2826, -687, 3078, 652, -3316, -645, 3562, 
634, -3796, -621, 4036, 630, -4251, -640, 4466, 648, 
-4667, -680, 4860, 695, -5028, -730, 5200, 778, -5342, 
-807, 5486, 866, -5600, -903, 5709, 957, -5788, -1011, 
5860, 1057, -5903, -1099, 5924, 1163, -5943, -1206, 5928, 
1243, -5894, -1275, 5849, 1316, -5767, -1332, 5678, 1350, 
-5565, -1359, 5435, 1367, -5292, -1354, 5113, 1334, -4930, 
-1305, 4724, 1261, -4511, -1216, 4278, 1148, -4023, -1069, 
3769, 985, -3486, -885, 3200, 780, -2902, -656, 2609, 
537, -2297, -381, 1971, 227, -1661, -74, 1336, -93, 
-1018, 272, 684, -467, -367, 650, 60, -853, 252, 
1051, -566, -1270, 859, 1472, -1150, -1683, 1429, 1891, 
-1690, -2091, 1948, 2290, -2183, -2492, 2423, 2685, -2629, 
-2874, 2826, 3053, -2991, -3230, 3158, 3395, -3304, -3541, 
3429, 3672, -3528, -3798, 3613, 3908, -3681, -4007, 3721, 
4087, -3758, -4149, 3773, 4184, -3761, -4212, 3740, 4225, 
-3691, -4224, 3634, 4197, -3562, -4161, 3477, 4095, -3365, 
-4014, 3256, 3929, -3137, -3813, 2985, 3683, -2839, -3534, 
2687, 3371, -2531, -3197, 2362, 3010, -2190, -2819, 2004, 
2602, -1829, -2390, 1637, 2158, -1459, -1918, 1281, 1669, 
-1089, -1421, 916, 1166, -746, -912, 567, 654, -413, 
-386, 260, 132, -105, 124, -47, -380, 175, 620, 
-295, -862, 419, 1093, -530, -1316, 623, 1531, -705, 
-1723, 789, 1913, -853, -2089, 911, 2254, -958, -2398, 
981, 2533, -1010, -2635, 1024, 2741, -1032, -2824, 1030, 
2879, -1025, -2930, 996, 2951, -977, -2977, 949, 2963, 
-897, -2931, 849, 2890, -796, -2835, 741, 2758, -685, 
-2654, 622, 2543, -554, -2418, 487, 2282, -416, -2116, 
331, 1952, -259, -1766, 189, 1562, -116, -1366, 36, 
1142, 31, -908, -110, 678, 168, -433, -250, 176, 
304, 80, -364, -338, 423, 602, -483, -867, 534, 
1147, -583, -1415, 629, 1687, -671, -1953, 696, 2224, 
-724, -2492, 757, 2767, -781, -3013, 787, 3271, -807, 
-3527, 816, 3769, -812, -4009, 819, 4233, -816, -4451, 
797, 4658, -795, -4862, 769, 5062, -753, -5241, 718, 
5407, -687, -5576, 657, 5718, -609, -5860, 565, 5986, 
-524, -6097, 465, 6205, -407, -6288, 341, 6373, -267, 
-6426, 199, 6476, -127, -6523, 54, 6553, 41, -6573, 
-119, 6571, 227, -6556, -316, 6545, 416, -6517, -520, 
6469, 625, -6404, -749, 6351, 864, -6274, -988, 6185, 
1102, -6081, -1233, 5979, 1364, -5857, -1487, 5741, 1620, 
-5602, -1752, 5450, 1887, -5314, -2031, 5147, 2169, -4986, 
-2299, 4808, 2439, -4635, -2579, 4463, 2697, -4264, -2841, 
4088, 2962, -3893, -3086, 3690, 3211, -3493, -3324, 3283, 
3426, -3086, -3523, 2875, 3628, -2675, -3714, 2467, 3807, 
-2264, -3871, 2059, 3945, -1855, -3999, 1656, 4034, -1456, 
-4069, 1259, 4094, -1062, -4114, 874, 4118, -699, -4100, 
521, 4089, -346, -4055, 165, 4003, -11, -3953, -159, 
3882, 298, -3804, -459, 3706, 595, -3611, -736, 3488, 
856, -3370, -985, 3244, 1114, -3098, -1217, 2947, 1330, 
-2779, -1424, 2613, 1529, -2435, -1625, 2262, 1715, -2071, 
-1789, 1889, 1878, -1691, -1950, 1495, 2016, -1295, -2090, 
1108, 2167, -910, -2220, 708, 2299, -524, -2358, 339, 
2423, -141, -2470, -34, 2542, 209, -2595, -360, 2670, 
526, -2733, -676, 2799, 814, -2865, -952, 2938, 1070, 
-3009, -1173, 3080, 1279, -3152, -1356, 3226, 1431, -3306, 
-1498, 3385, 1545, -3474, -1576, 3572, 1608, -3651, -1623, 
3754, 1613, -3844, -1605, 3942, 1573, -4037, -1537, 4130, 
1492, -4227, -1434, 4329, 1365, -4422, -1288, 4507, 1195, 
-4609, -1095, 4701, 1007, -4782, -880, 4859, 770, -4942, 
-641, 5014, 528, -5069, -397, 5129, 255, -5167, -122, 
5219, -12, -5240, 166, 5267, -295, -5266, 435, 5262, 
-583, -5260, 709, 5230, -847, -5187, 981, 5123, -1098, 
-5059, 1225, 4987, -1347, -4880, 1469, 4773, -1579, -4642, 
1674, 4500, -1779, -4346, 1860, 4173, -1949, -3984, 2035, 
3783, -2110, -3566, 2173, 3341, -2246, -3097, 2296, 2833, 
-2339, -2574, 2392, 2289, -2430, -2002, 2468, 1696, -2498, 
-1395, 2518, 1089, -2539, -759, 2544, 438, -2559, -100, 
2559, -234, -2560, 577, 2557, -916, -2540, 1245, 2525, 
-1582, -2519, 1910, 2498, -2236, -2460, 2574, 2440, -2885, 
-2416, 3203, 2373, -3504, -2338, 3787, 2292, -4070, -2244, 
4336, 2188, -4590, -2129, 4825, 2071, -5061, -1997, 5277, 
1938, -5464, -1861, 5652, 1777, -5811, -1685, 5956, 1590, 
-6077, -1496, 6185, 1391, -6273, -1283, 6341, 1159, -6406, 
-1033, 6438, 896, -6454, -757, 6443, 611, -6428, -461, 
6393, 305, -6337, -128, 6273, -47, -6183, 217, 6084, 
-406, -5973, 603, 5848, -794, -5708, 996, 5546, -1196, 
-5397, 1396, 5220, -1615, -5039, 1830, 4842, -2045, -4659, 
2251, 4454, -2453, -4244, 2677, 4041, -2877, -3827, 3077, 
3623, -3273, -3401, 3462, 3191, -3656, -2979, 3822, 2769, 
-3994, -2565, 4152, 2362, -4284, -2156, 4417, 1959, -4540, 
-1779, 4642, 1599, -4722, -1419, 4782, 1245, -4839, -1089, 
4870, 935, -4895, -778, 4888, 648, -4852, -518, 4813, 
404, -4746, -289, 4669, 189, -4570, -90, 4444, 3, 
-4301, 80, 4131, -145, -3951, 201, 3765, -258, -3552, 
301, 3319, -340, -3068, 366, 2805, -390, -2548, 409, 
2264, -425, -1976, 426, 1677, -433, -1375, 423, 1063, 
-412, -756, 414, 432, -389, -127, 375, -170, -354, 
479, 327, -777, -314, 1056, 287, -1335, -252, 1590, 
215, -1830, -192, 2070, 165, -2273, -132, 2474, 96, 
-2644, -69, 2793, 42, -2922, -10, 3021, -32, -3091, 
55, 3139, -85, -3168, 128, 3160, -143, -3129, 183, 
3068, -204, -2991, 242, 2876, -276, -2730, 303, 2558, 
-336, -2370, 368, 2161, -396, -1926, 415, 1666, -462, 
-1376, 487, 1079, -514, -767, 559, 427, -599, -86, 
626, -270, -661, 636, 702, -1020, -759, 1399, 804, 
-1772, -850, 2166, 893, -2534, -941, 2916, 1000, -3290, 
-1053, 3646, 1111, -3984, -1165, 4331, 1233, -4641, -1303, 
4946, 1363, -5238, -1430, 5497, 1501, -5722, -1580, 5951, 
1655, -6127, -1729, 6299, 1805, -6430, -1892, 6525, 1983, 
-6603, -2067, 6635, 2143, -6653, -2237, 6637, 2318, -6582, 
-2400, 6501, 2495, -6380, -2571, 6244, 2651, -6056, -2751, 
5867, 2828, -5627, -2915, 5365, 2994, -5086, -3071, 4786, 
3136, -4454, -3216, 4100, 3295, -3732, -3355, 3343, 3419, 
-2935, -3471, 2518, 3524, -2100, -3587, 1668, 3626, -1216, 
-3672, 766, 3703, -324, -3729, -134, 3756, 576, -3770, 
-1031, 3776, 1476, -3777, -1908, 3771, 2331, -3753, -2748, 
3727, 3147, -3691, -3531, 3664, 3910, -3612, -4264, 3551, 
4594, -3495, -4907, 3426, 5204, -3348, -5480, 3253, 5726, 
-3161, -5963, 3051, 6165, -2923, -6356, 2807, 6503, -2676, 
-6642, 2532, 6755, -2398, -6850, 2237, 6912, -2075, -6961, 
1918, 6980, -1739, -6974, 1557, 6951, -1381, -6914, 1192, 
6856, -1002, -6768, 801, 6665, -608, -6567, 404, 6437, 
-200, -6290, 10, 6139, 197, -5970, -399, 5791, 600, 
-5599, -798, 5410, 990, -5202, -1173, 4993, 1358, -4783, 
-1535, 4568, 1711, -4340, -1887, 4123, 2038, -3901, -2193, 
3682, 2334, -3459, -2458, 3224, 2585, -3019, -2698, 2790, 
2788, -2577, -2885, 2378, 2954, -2164, -3015, 1972, 3073, 
-1772, -3110, 1577, 3137, -1405, -3143, 1222, 3145, -1045, 
-3142, 882, 3114, -717, -3079, 565, 3023, -425, -2957, 
290, 2885, -154, -2800, 30, 2708, 85, -2596, -197, 
2474, 302, -2366, -400, 2230, 495, -2089, -582, 1951, 
659, -1809, -725, 1642, 792, -1502, -853, 1338, 902, 
-1178, -943, 1034, 981, -876, -998, 719, 1028, -573, 
-1036, 421, 1045, -280, -1037, 159, 1034, -31, -1019, 
-87, 996, 199, -965, -289, 922, 369, -873, -455, 
826, 515, -751, -559, 682, 593, -604, -614, 512, 
634, -427, -628, 328, 616, -206, -583, 101, 529, 
35, -472, -163, 403, 290, -320, -437, 215, 592, 
-116, -740, -12, 903, 133, -1066, -277, 1228, 418, 
-1387, -571, 1558, 739, -1726, -911, 1900, 1085, -2068, 
-1253, 2235, 1425, -2403, -1614, 2555, 1781, -2729, -1962, 
2870, 2136, -3022, -2305, 3175, 2457, -3309, -2613, 3438, 
2762, -3558, -2911, 3667, 3031, -3771, -3158, 3853, 3260, 
-3932, -3348, 4015, 3422, -4059, -3499, 4102, 3546, -4130, 
-3577, 4158, 3598, -4155, -3592, 4151, 3576, -4130, -3552, 
4088, 3494, -4049, -3441, 3984, 3351, -3899, -3251, 3816, 
3135, -3712, -3012, 3612, 2868, -3483, -2713, 3354, 2547, 
-3211, -2363, 3050, 2176, -2897, -1971, 2733, 1750, -2557, 
-1537, 2379, 1316, -2180, -1074, 1996, 838, -1798, -610, 
1616, 364, -1410, -128, 1217, -108, -1038, 326, 841, 
-553, -646, 780, 465, -988, -286, 1195, 110, -1395, 
53, 1584, -218, -1750, 372, 1906, -527, -2056, 661, 
2181, -788, -2298, 909, 2383, -1023, -2475, 1127, 2530, 
-1222, -2569, 1301, 2599, -1369, -2614, 1425, 2594, -1477, 
-2566, 1513, 2523, -1553, -2443, 1577, 2367, -1593, -2271, 
1595, 2148, -1597, -2015, 1571, 1858, -1569, -1698, 1539, 
1528, -1502, -1335, 1480, 1126, -1437, -925, 1387, 705, 
-1340, -478, 1288, 242, -1232, 5, 1170, -241, -1119, 
487, 1057, -733, -1006, 982, 946, -1222, -880, 1464, 
817, -1692, -760, 1922, 702, -2153, -652, 2363, 595, 
-2571, -541, 2752, 486, -2935, -431, 3119, 375, -3270, 
-332, 3417, 282, -3530, -231, 3655, 191, -3744, -136, 
3831, 93, -3897, -32, 3932, -17, -3960, 66, 3979, 
-118, -3978, 171, 3953, -216, -3905, 287, 3854, -344, 
-3784, 406, 3703, -469, -3602, 549, 3493, -615, -3363, 
693, 3222, -774, -3064, 858, 2911, -953, -2741, 1047, 
2560, -1132, -2362, 1238, 2169, -1342, -1964, 1448, 1764, 
-1553, -1548, 1657, 1347, -1748, -1136, 1854, 922, -1969, 
-711, 2062, 515, -2172, -318, 2260, 118, -2357, 75, 
2432, -248, -2524, 427, 2600, -600, -2661, 750, 2705, 
-891, -2759, 1027, 2793, -1146, -2811, 1266, 2828, -1359, 
-2821, 1445, 2792, -1495, -2773, 1564, 2718, -1596, -2656, 
1616, 2571, -1622, -2465, 1619, 2339, -1584, -2203, 1553, 
2062, -1489, -1885, 1426, 1692, -1334, -1481, 1251, 1257, 
-1131, -1023, 1017, 761, -880, -500, 728, 209, -565, 
81, 386, -404, -213, 719, 30, -1045, 163, 1384, 
-376, -1738, 582, 2091, -796, -2445, 1008, 2794, -1227, 
-3141, 1463, 3497, -1672, -3845, 1905, 4185, -2127, -4527, 
2344, 4846, -2566, -5163, 2781, 5469, -2984, -5747, 3186, 
6024, -3381, -6271, 3561, 6497, -3733, -6713, 3910, 6894, 
-4067, -7055, 4210, 7183, -4330, -7298, 4454, 7390, -4567, 
-7446, 4664, 7469, -4737, -7475, 4802, 7440, -4858, -7387, 
4892, 7299, -4912, -7185, 4910, 7037, -4899, -6862, 4870, 
6665, -4827, -6448, 4773, 6197, -4694, -5926, 4602, 5631, 
-4507, -5319, 4383, 4994, -4265, -4645, 4111, 4276, -3963, 
-3911, 3801, 3520, -3624, -3134, 3429, 2721, -3247, -2317, 
3041, 1917, -2822, -1516, 2596, 1112, -2384, -708, 2149, 
321, -1919, 70, 1672, -430, -1440, 800, 1200, -1140, 
-966, 1457, 721, -1766, -475, 2049, 251, -2315, -16, 
2545, -205, -2764, 439, 2951, -652, -3105, 849, 3247, 
-1055, -3347, 1247, 3417, -1441, -3469, 1622, 3488, -1783, 
-3467, 1941, 3432, -2090, -3366, 2218, 3275, -2346, -3145, 
2466, 2995, -2561, -2818, 2657, 2636, -2737, -2412, 2806, 
2167, -2880, -1911, 2929, 1648, -2956, -1350, 2988, 1056, 
-3019, -733, 3022, 407, -3028, -84, 3018, -257, -3002, 
598, 2984, -940, -2951, 1276, 2927, -1625, -2876, 1960, 
2836, -2289, -2797, 2611, 2736, -2917, -2689, 3214, 2630, 
-3510, -2568, 3784, 2495, -4025, -2448, 4279, 2386, -4492, 
-2313, 4704, 2253, -4888, -2198, 5043, 2137, -5184, -2067, 
5315, 2022, -5413, -1968, 5487, 1909, -5537, -1867, 5578, 
1824, -5599, -1778, 5595, 1731, -5564, -1692, 5527, 1666, 
-5460, -1634, 5392, 1589, -5300, -1566, 5192, 1546, -5055, 
-1521, 4926, 1490, -4783, -1467, 4631, 1459, -4461, -1430, 
4280, 1419, -4113, -1407, 3924, 1389, -3741, -1371, 3566, 
1354, -3370, -1335, 3186, 1324, -3003, -1304, 2837, 1286, 
-2668, -1271, 2498, 1251, -2339, -1237, 2179, 1210, -2043, 
-1203, 1910, 1170, -1786, -1164, 1674, 1141, -1562, -1125, 
1483, 1093, -1406, -1077, 1335, 1070, -1281, -1058, 1237, 
1042, -1208, -1036, 1185, 1033, -1164, -1023, 1174, 1031, 
-1181, -1047, 1201, 1048, -1228, -1078, 1266, 1095, -1315, 
-1141, 1371, 1170, -1426, -1227, 1488, 1284, -1549, -1357, 
1621, 1434, -1688, -1524, 1764, 1613, -1830, -1721, 1913, 
1845, -1974, -1971, 2046, 2113, -2103, -2270, 2174, 2415, 
-2229, -2589, 2270, 2777, -2327, -2967, 2361, 3161, -2403, 
-3368, 2414, 3575, -2434, -3806, 2451, 4031, -2452, -4248, 
2436, 4493, -2431, -4727, 2410, 4978, -2367, -5210, 2330, 
5458, -2282, -5688, 2231, 5920, -2162, -6163, 2090, 6389, 
-2016, -6600, 1927, 6816, -1831, -7022, 1735, 7215, -1641, 
-7396, 1530, 7556, -1423, -7711, 1308, 7844, -1194, -7964, 
1067, 8065, -951, -8151, 822, 8210, -688, -8256, 565, 
8271, -436, -8273, 324, 8254, -185, -8211, 62, 8150, 
63, -8070, -180, 7963, 302, -7831, -417, 7672, 533, 
-7508, -649, 7314, 766, -7108, -866, 6876, 971, -6625, 
-1075, 6370, 1181, -6093, -1294, 5800, 1383, -5494, -1481, 
5189, 1592, -4858, -1685, 4529, 1778, -4193, -1877, 3849, 
1975, -3496, -2075, 3149, 2168, -2815, -2268, 2458, 2366, 
-2123, -2465, 1796, 2565, -1470, -2675, 1136, 2782, -843, 
-2885, 533, 2992, -246, -3110, -23, 3220, 271, -3340, 
-517, 3459, 740, -3581, -949, 3710, 1136, -3835, -1304, 
3962, 1454, -4080, -1585, 4217, 1699, -4347, -1807, 4480, 
1882, -4613, -1949, 4732, 1978, -4868, -2014, 4982, 2021, 
-5109, -2012, 5225, 2005, -5345, -1964, 5459, 1934, -5559, 
-1876, 5661, 1821, -5759, -1750, 5841, 1675, -5917, -1591, 
5982, 1506, -6040, -1430, 6089, 1349, -6129, -1273, 6155, 
1196, -6170, -1124, 6159, 1046, -6149, -991, 6128, 935, 
-6099, -896, 6035, 879, -5978, -859, 5892, 852, -5811, 
-852, 5692, 884, -5583, -911, 5448, 966, -5289, -1029, 
5133, 1122, -4968, -1221, 4775, 1333, -4582, -1451, 4370, 
1589, -4159, -1746, 3933, 1909, -3699, -2073, 3447, 2259, 
-3205, -2454, 2949, 2667, -2690, -2865, 2433, 3088, -2161, 
-3305, 1903, 3520, -1628, -3730, 1357, 3955, -1096, -4159, 
843, 4381, -589, -4576, 337, 4767, -91, -4952, -144, 
5136, 388, -5288, -595, 5445, 816, -5571, -1011, 5687, 
1205, -5788, -1379, 5867, 1537, -5915, -1677, 5952, 1827, 
-5976, -1934, 5982, 2048, -5948, -2143, 5910, 2215, -5840, 
-2282, 5751, 2322, -5629, -2358, 5504, 2367, -5353, -2374, 
5179, 2375, -5000, -2352, 4781, 2308, -4559, -2257, 4322, 
2203, -4074, -2129, 3814, 2041, -3540, -1965, 3244, 1857, 
-2960, -1753, 2656, 1650, -2364, -1527, 2063, 1396, -1760, 
-1282, 1458, 1160, -1166, -1031, 867, 888, -582, -764, 
309, 642, -35, -507, -206, 395, 452, -272, -680, 
176, 886, -66, -1078, -41, 1260, 124, -1411, -199, 
1554, 282, -1676, -351, 1758, 399, -1843, -446, 1902, 
488, -1936, -501, 1949, 516, -1929, -529, 1905, 517, 
-1863, -493, 1796, 472, -1706, -442, 1600, 395, -1488, 
-323, 1364, 271, -1217, -183, 1053, 112, -892, -22, 
710, -76, -529, 185, 326, -291, -125, 412, -60, 
-527, 269, 653, -471, -771, 674, 897, -873, -1018, 
1071, 1148, -1259, -1284, 1437, 1405, -1610, -1525, 1776, 
1646, -1929, -1775, 2064, 1883, -2196, -1987, 2309, 2100, 
-2420, -2188, 2509, 2286, -2582, -2369, 2645, 2450, -2687, 
-2533, 2722, 2593, -2732, -2644, 2737, 2699, -2723, -2729, 
2681, 2768, -2649, -2789, 2591, 2790, -2529, -2797, 2446, 
2790, -2350, -2781, 2255, 2755, -2146, -2711, 2035, 2670, 
-1919, -2629, 1776, 2556, -1646, -2488, 1512, 2423, -1378, 
-2343, 1239, 2248, -1096, -2149, 961, 2039, -830, -1934, 
693, 1804, -571, -1685, 445, 1554, -323, -1425, 215, 
1281, -102, -1138, 5, 972, 67, -825, -153, 669, 
228, -504, -270, 325, 325, -167, -367, -14, 384, 
188, -399, -369, 416, 541, -398, -737, 395, 911, 
-363, -1101, 321, 1294, -286, -1480, 228, 1659, -168, 
-1851, 95, 2039, -18, -2234, -69, 2413, 162, -2607, 
-276, 2787, 383, -2956, -481, 3148, 601, -3327, -728, 
3498, 850, -3655, -971, 3829, 1100, -3980, -1230, 4141, 
1372, -4283, -1498, 4437, 1632, -4573, -1766, 4684, 1904, 
-4818, -2021, 4928, 2161, -5024, -2293, 5113, 2412, -5192, 
-2535, 5249, 2670, -5313, -2786, 5351, 2913, -5386, -3017, 
5398, 3138, -5406, -3251, 5403, 3359, -5376, -3452, 5335, 
3558, -5273, -3661, 5193, 3739, -5116, -3830, 5004, 3912, 
-4887, -4009, 4748, 4082, -4604, -4156, 4430, 4219, -4246, 
-4284, 4050, 4334, -3841, -4393, 3613, 4437, -3373, -4470, 
3103, 4517, -2836, -4544, 2567, 4567, -2278, -4569, 1986, 
4583, -1665, -4581, 1363, 4572, -1037, -4550, 718, 4522, 
-383, -4472, 48, 4422, 271, -4378, -616, 4302, 943, 
-4224, -1273, 4130, 1586, -4021, -1901, 3906, 2215, -3785, 
-2516, 3649, 2797, -3501, -3067, 3334, 3340, -3168, -3588, 
2990, 3818, -2793, -4028, 2589, 4220, -2358, -4398, 2145, 
4559, -1905, -4691, 1654, 4818, -1409, -4904, 1144, 4971, 
-891, -5017, 614, 5046, -339, -5051, 60, 5020, 224, 
-4977, -512, 4901, 797, -4815, -1065, 4706, 1353, -4566, 
-1623, 4406, 1902, -4230, -2154, 4036, 2420, -3829, -2657, 
3592, 2902, -3357, -3117, 3096, 3330, -2829, -3520, 2551, 
3702, -2254, -3878, 1958, 4014, -1652, -4155, 1353, 4264, 
-1045, -4340, 728, 4420, -432, -4464, 121, 4495, 175, 
-4494, -462, 4470, 758, -4424, -1031, 4360, 1288, -4288, 
-1530, 4179, 1767, -4039, -1987, 3893, 2193, -3723, -2383, 
3520, 2543, -3314, -2694, 3081, 2824, -2827, -2920, 2567, 
3012, -2288, -3076, 1997, 3113, -1696, -3134, 1367, 3128, 
-1052, -3111, 723, 3059, -381, -2999, 34, 2909, 313, 
-2815, -663, 2678, 1019, -2548, -1364, 2383, 1716, -2223, 
-2059, 2033, 2380, -1839, -2722, 1629, 3041, -1413, -3351, 
1182, 3644, -960, -3928, 727, 4202, -485, -4463, 230, 
4708, 4, -4932, -250, 5150, 491, -5337, -719, 5531, 
964, -5690, -1181, 5834, 1400, -5963, -1604, 6079, 1811, 
-6167, -1995, 6245, 2161, -6306, -2324, 6351, 2488, -6378, 
-2614, 6391, 2739, -6389, -2856, 6371, 2948, -6346, -3027, 
6294, 3086, -6249, -3147, 6190, 3181, -6114, -3191, 6026, 
3210, -5939, -3200, 5852, 3193, -5756, -3171, 5649, 3121, 
-5535, -3081, 5424, 3025, -5302, -2956, 5178, 2899, -5049, 
-2822, 4929, 2735, -4804, -2656, 4688, 2566, -4555, -2477, 
4426, 2373, -4305, -2293, 4183, 2206, -4069, -2106, 3953, 
2026, -3825, -1949, 3712, 1873, -3597, -1808, 3475, 1742, 
-3360, -1679, 3234, 1615, -3130, -1580, 3014, 1535, -2891, 
-1495, 2778, 1479, -2645, -1458, 2540, 1441, -2413, -1447, 
2289, 1439, -2163, -1455, 2030, 1477, -1898, -1492, 1759, 
1520, -1621, -1549, 1464, 1569, -1318, -1608, 1169, 1640, 
-1018, -1687, 858, 1723, -692, -1757, 535, 1810, -366, 
-1840, 206, 1877, -29, -1909, -134, 1940, 309, -1964, 
-473, 1967, 651, -1983, -824, 2005, 986, -2005, -1152, 
1992, 1305, -1975, -1473, 1963, 1612, -1941, -1759, 1911, 
1902, -1863, -2027, 1829, 2159, -1778, -2266, 1718, 2373, 
-1664, -2455, 1597, 2550, -1519, -2613, 1443, 2672, -1372, 
-2707, 1284, 2751, -1217, -2761, 1120, 2774, -1046, -2761, 
971, 2744, -891, -2715, 823, 2664, -746, -2608, 682, 
2526, -635, -2444, 581, 2356, -545, -2252, 511, 2138, 
-490, -2012, 474, 1886, -456, -1744, 479, 1590, -491, 
-1450, 518, 1294, -574, -1137, 625, 979, -684, -828, 
765, 657, -863, -516, 969, 360, -1092, -213, 1218, 
66, -1347, 70, 1492, -196, -1650, 310, 1811, -435, 
-1984, 524, 2156, -628, -2348, 693, 2523, -766, -2723, 
825, 2911, -861, -3099, 896, 3278, -914, -3456, 915, 
3646, -910, -3812, 887, 3982, -857, -4133, 806, 4271, 
-752, -4416, 686, 4537, -610, -4656, 521, 4744, -428, 
-4829, 331, 4889, -233, -4941, 115, 4972, 0, -4987, 
-121, 4984, 227, -4956, -351, 4907, 466, -4858, -588, 
4779, 692, -4684, -804, 4567, 913, -4438, -1004, 4289, 
1101, -4116, -1180, 3940, 1244, -3753, -1318, 3560, 1377, 
-3345, -1413, 3118, 1442, -2885, -1471, 2650, 1471, -2398, 
-1472, 2158, 1458, -1908, -1439, 1663, 1403, -1414, -1341, 
1156, 1299, -929, -1219, 693, 1149, -450, -1067, 231, 
987, -23, -882, -167, 782, 355, -684, -525, 574, 
678, -450, -817, 345, 951, -239, -1048, 128, 1142, 
-21, -1205, -84, 1264, 175, -1288, -275, 1317, 348, 
-1306, -436, 1283, 496, -1244, -554, 1195, 597, -1133, 
-638, 1034, 668, -934, -670, 831, 686, -711, -677, 
580, 654, -423, -620, 278, 577, -122, -514, -41, 
452, 204, -368, -373, 288, 536, -187, -707, 89, 
862, 22, -1023, -135, 1176, 248, -1320, -368, 1442, 
488, -1566, -603, 1678, 730, -1786, -847, 1870, 966, 
-1939, -1087, 1996, 1193, -2039, -1289, 2075, 1369, -2081, 
-1456, 2082, 1526, -2067, -1585, 2030, 1634, -1976, -1651, 
1907, 1671, -1823, -1681, 1725, 1681, -1624, -1653, 1504, 
1620, -1374, -1565, 1226, 1491, -1080, -1412, 915, 1323, 
-751, -1222, 581, 1109, -421, -975, 241, 845, -77, 
-702, -97, 554, 257, -391, -421, 232, 571, -75, 
-714, -101, 842, 251, -975, -417, 1091, 575, -1182, 
-712, 1273, 856, -1350, -986, 1408, 1115, -1437, -1220, 
1469, 1318, -1475, -1391, 1464, 1457, -1429, -1491, 1389, 
1519, -1332, -1523, 1250, 1504, -1159, -1466, 1046, 1413, 
-914, -1322, 773, 1220, -631, -1108, 469, 956, -302, 
-797, 126, 615, 64, -403, -260, 197, 448, 46, 
-639, -291, 837, 556, -1032, -834, 1216, 1114, -1398, 
-1396, 1559, 1690, -1726, -1990, 1875, 2276, -2014, -2582, 
2148, 2870, -2247, -3150, 2337, 3426, -2413, -3688, 2467, 
3930, -2497, -4173, 2513, 4388, -2499, -4584, 2463, 4753, 
-2400, -4905, 2320, 5021, -2212, -5116, 2083, 5187, -1919, 
-5237, 1757, 5243, -1547, -5225, 1340, 5188, -1103, -5101, 
844, 4989, -568, -4862, 276, 4694, 25, -4493, -350, 
4284, 674, -4035, -1009, 3767, 1340, -3473, -1699, 3151, 
2046, -2834, -2397, 2485, 2729, -2138, -3084, 1761, 3404, 
-1387, -3729, 1010, 4056, -641, -4353, 269, 4628, 105, 
-4887, -459, 5135, 809, -5362, -1161, 5565, 1480, -5728, 
-1770, 5878, 2055, -6004, -2302, 6083, 2517, -6152, -2714, 
6178, 2886, -6171, -3012, 6125, 3105, -6070, -3160, 5966, 
3188, -5825, -3169, 5668, 3113, -5470, -3015, 5246, 2893, 
-4995, -2719, 4705, 2499, -4400, -2267, 4052, 1992, -3705, 
-1679, 3312, 1322, -2913, -958, 2498, 554, -2059, -132, 
1608, -313, -1134, 768, 662, -1240, -192, 1733, -300, 
-2237, 778, 2745, -1280, -3247, 1753, 3742, -2235, -4229, 
2707, 4715, -3174, -5194, 3617, 5647, -4050, -6084, 4465, 
6499, -4867, -6881, 5241, 7234, -5597, -7552, 5933, 7842, 
-6237, -8081, 6517, 8293, -6769, -8457, 6994, 8594, -7193, 
-8674, 7356, 8696, -7493, -8700, 7595, 8643, -7663, -8539, 
7699, 8398, -7711, -8202, 7687, 7974, -7643, -7703, 7563, 
7392, -7453, -7027, 7309, 6640, -7155, -6229, 6967, 5773, 
-6758, -5294, 6516, 4804, -6276, -4282, 6001, 3745, -5710, 
-3192, 5414, 2633, -5095, -2059, 4775, 1493, -4431, -924, 
4086, 371, -3755, 179, 3392, -719, -3048, 1222, 2696, 
-1721, -2362, 2199, 2023, -2641, -1684, 3051, 1357, -3420, 
-1040, 3759, 750, -4070, -452, 4334, 177, -4556, 64, 
4731, -304, -4869, 533, 4945, -722, -4985, 901, 4990, 
-1060, -4942, 1201, 4841, -1314, -4697, 1402, 4527, -1473, 
-4304, 1515, 4034, -1537, -3731, 1531, 3401, -1496, -3039, 
1452, 2633, -1386, -2213, 1293, 1769, -1171, -1306, 1047, 
824, -892, -322, 721, -182, -526, 695, 332, -1208, 
-98, 1712, -122, -2224, 370, 2722, -620, -3203, 884, 
3666, -1163, -4129, 1452, 4552, -1723, -4946, 2022, 5331, 
-2307, -5681, 2605, 5996, -2894, -6270, 3175, 6510, -3451, 
-6719, 3733, 6890, -4000, -7028, 4278, 7122, -4531, -7176, 
4773, 7188, -5006, -7169, 5220, 7096, -5418, -7001, 5615, 
6859, -5778, -6693, 5943, 6489, -6079, -6256, 6201, 5986, 
-6294, -5699, 6388, 5378, -6442, -5046, 6487, 4677, -6507, 
-4304, 6503, 3921, -6493, -3520, 6453, 3126, -6392, -2712, 
6306, 2292, -6201, -1891, 6083, 1487, -5952, -1085, 5783, 
701, -5617, -308, 5426, -52, -5217, 398, 4997, -723, 
-4756, 1033, 4499, -1332, -4244, 1602, 3972, -1844, -3694, 
2047, 3398, -2238, -3096, 2413, 2799, -2547, -2488, 2668, 
2170, -2745, -1862, 2809, 1558, -2833, -1235, 2850, 931, 
-2830, -625, 2788, 331, -2738, -28, 2658, -257, -2550, 
522, 2445, -797, -2303, 1045, 2168, -1278, -2015, 1513, 
1842, -1715, -1667, 1910, 1490, -2092, -1315, 2257, 1135, 
-2398, -943, 2527, 768, -2638, -588, 2711, 408, -2787, 
-229, 2831, 69, -2862, 73, 2873, -213, -2853, 359, 
2829, -473, -2778, 586, 2701, -684, -2627, 780, 2528, 
-849, -2406, 907, 2268, -964, -2116, 1011, 1953, -1038, 
-1775, 1049, 1597, -1071, -1398, 1069, 1206, -1061, -989, 
1048, 772, -1041, -546, 1014, 326, -1010, -109, 985, 
-122, -970, 345, 955, -552, -931, 767, 930, -979, 
-926, 1178, 945, -1380, -951, 1557, 982, -1730, -1027, 
1888, 1069, -2040, -1138, 2162, 1200, -2277, -1302, 2391, 
1405, -2463, -1518, 2536, 1643, -2591, -1792, 2623, 1941, 
-2635, -2111, 2643, 2296, -2607, -2485, 2585, 2701, -2521, 
-2914, 2457, 3127, -2360, -3359, 2254, 3583, -2141, -3812, 
1998, 4055, -1849, -4289, 1690, 4525, -1522, -4754, 1343, 
4972, -1150, -5182, 944, 5388, -745, -5569, 539, 5751, 
-309, -5908, 103, 6050, 113, -6172, -339, 6271, 547, 
-6359, -766, 6411, 968, -6441, -1178, 6443, 1377, -6418, 
-1557, 6365, 1736, -6287, -1911, 6174, 2054, -6043, -2214, 
5873, 2341, -5685, -2459, 5458, 2558, -5215, -2658, 4941, 
2729, -4648, -2779, 4320, 2833, -3972, -2852, 3610, 2876, 
-3212, -2881, 2810, 2857, -2395, -2823, 1962, 2792, -1515, 
-2722, 1053, 2651, -596, -2583, 134, 2479, 341, -2381, 
-799, 2273, 1273, -2154, -1720, 2021, 2183, -1892, -2619, 
1764, 3048, -1618, -3460, 1475, 3860, -1333, -4243, 1183, 
4599, -1038, -4935, 896, 5253, -758, -5547, 628, 5804, 
-495, -6040, 367, 6257, -242, -6435, 134, 6577, -39, 
-6708, -63, 6807, 143, -6876, -227, 6916, 283, -6926, 
-355, 6894, 403, -6862, -435, 6798, 465, -6699, -494, 
6580, 491, -6447, -510, 6287, 497, -6125, -478, 5932, 
465, -5730, -446, 5514, 408, -5275, -371, 5045, 338, 
-4794, -296, 4553, 248, -4303, -196, 4044, 154, -3797, 
-107, 3539, 73, -3290, -29, 3051, 2, -2823, 30, 
2593, -54, -2381, 89, 2182, -97, -1991, 96, 1804, 
-103, -1636, 94, 1485, -70, -1347, 44, 1222, -5, 
-1118, -39, 1023, 92, -936, -147, 868, 218, -818, 
-303, 769, 389, -749, -497, 739, 600, -732, -707, 
735, 829, -744, -955, 758, 1087, -787, -1202, 827, 
1346, -856, -1485, 899, 1616, -943, -1739, 981, 1870, 
-1022, -2013, 1068, 2132, -1101, -2241, 1132, 2358, -1157, 
-2464, 1177, 2558, -1200, -2645, 1202, 2727, -1211, -2789, 
1197, 2846, -1190, -2888, 1163, 2912, -1135, -2910, 1093, 
2920, -1048, -2904, 990, 2869, -915, -2812, 838, 2758, 
-760, -2670, 668, 2568, -563, -2469, 469, 2341, -359, 
-2207, 249, 2042, -126, -1893, 16, 1710, 98, -1524, 
-218, 1320, 345, -1124, -460, 903, 575, -687, -675, 
463, 795, -216, -892, -4, 980, 238, -1071, -483, 
1149, 716, -1228, -953, 1295, 1169, -1355, -1400, 1398, 
1619, -1430, -1822, 1465, 2031, -1484, -2213, 1503, 2391, 
-1503, -2571, 1483, 2725, -1470, -2864, 1455, 2994, -1432, 
-3117, 1393, 3218, -1353, -3287, 1307, 3369, -1254, -3427, 
1204, 3465, -1146, -3486, 1100, 3493, -1041, -3479, 988, 
3464, -950, -3424, 889, 3378, -855, -3317, 825, 3248, 
-798, -3166, 773, 3078, -762, -2976, 763, 2863, -788, 
-2744, 809, 2624, -841, -2500, 885, 2373, -938, -2232, 
1012, 2109, -1094, -1972, 1192, 1841, -1291, -1722, 1424, 
1592, -1551, -1468, 1686, 1356, -1850, -1240, 2003, 1130, 
-2182, -1040, 2354, 946, -2540, -867, 2737, 809, -2926, 
-746, 3137, 693, -3338, -656, 3530, 622, -3732, -589, 
3924, 588, -4110, -577, 4301, 582, -4472, -598, 4637, 
622, -4788, -647, 4927, 672, -5056, -728, 5166, 760, 
-5263, -813, 5339, 873, -5403, -925, 5441, 976, -5455, 
-1036, 5454, 1095, -5442, -1142, 5405, 1202, -5343, -1245, 
5260, 1286, -5144, -1336, 5028, 1368, -4873, -1399, 4723, 
1405, -4543, -1419, 4336, 1422, -4117, -1420, 3889, 1394, 
-3655, -1375, 3404, 1344, -3141, -1297, 2867, 1242, -2589, 
-1168, 2305, 1099, -2029, -1015, 1749, 918, -1462, -810, 
1194, 711, -920, -582, 666, 460, -405, -340, 174, 
195, 50, -58, -255, -73, 452, 223, -614, -360, 
770, 508, -890, -646, 1000, 781, -1071, -920, 1121, 
1041, -1157, -1172, 1154, 1289, -1136, -1400, 1069, 1487, 
-995, -1590, 899, 1655, -764, -1731, 603, 1778, -430, 
-1827, 224, 1853, -6, -1869, -242, 1864, 492, -1854, 
-769, 1821, 1054, -1774, -1360, 1711, 1667, -1638, -1984, 
1555, 2318, -1440, -2641, 1324, 2957, -1205, -3282, 1059, 
3605, -909, -3898, 744, 4196, -582, -4491, 391, 4749, 
-215, -5009, 16, 5237, 175, -5445, -377, 5626, 578, 
-5767, -792, 5906, 996, -6000, -1199, 6070, 1397, -6104, 
-1598, 6097, 1789, -6063, -1977, 5997, 2147, -5894, -2323, 
5758, 2481, -5584, -2624, 5382, 2763, -5136, -2892, 4862, 
3011, -4553, -3115, 4224, 3197, -3870, -3283, 3480, 3337, 
-3064, -3389, 2620, 3422, -2153, -3435, 1690, 3440, -1197, 
-3434, 696, 3416, -170, -3384, -340, 3349, 878, -3291, 
-1404, 3219, 1916, -3157, -2447, 3074, 2962, -2984, -3461, 
2884, 3945, -2797, -4423, 2682, 4878, -2578, -5307, 2468, 
5718, -2368, -6102, 2266, 6450, -2162, -6769, 2054, 7065, 
-1968, -7323, 1883, 7548, -1800, -7731, 1718, 7886, -1655, 
-7996, 1593, 8069, -1553, -8110, 1509, 8117, -1483, -8081, 
1474, 8000, -1468, -7897, 1468, 7745, -1496, -7569, 1522, 
7348, -1560, -7113, 1626, 6841, -1684, -6539, 1760, 6218, 
-1844, -5871, 1939, 5502, -2032, -5118, 2140, 4719, -2259, 
-4313, 2383, 3883, -2505, -3450, 2633, 3030, -2747, -2588, 
2874, 2154, -3006, -1734, 3139, 1305, -3245, -896, 3359, 
503, -3467, -112, 3577, -265, -3672, 616, 3742, -944, 
-3817, 1259, 3875, -1530, -3910, 1804, 3946, -2040, -3955, 
2240, 3950, -2422, -3920, 2575, 3894, -2683, -3838, 2788, 
3759, -2844, -3671, 2876, 3550, -2894, -3429, 2864, 3287, 
-2827, -3123, 2745, 2940, -2647, -2748, 2540, 2530, -2384, 
-2307, 2227, 2070, -2060, -1820, 1855, 1543, -1658, -1270, 
1434, 989, -1208, -715, 969, 408, -733, -119, 486, 
-184, -236, 471, 2, -782, 249, 1067, -480, -1354, 
703, 1641, -912, -1925, 1105, 2194, -1303, -2437, 1477, 
2685, -1616, -2921, 1759, 3133, -1877, -3326, 1968, 3509, 
-2045, -3664, 2099, 3794, -2125, -3920, 2113, 4012, -2102, 
-4092, 2050, 4151, -1994, -4181, 1889, 4182, -1777, -4177, 
1649, 4148, -1479, -4077, 1303, 4005, -1116, -3917, 898, 
3789, -664, -3659, 416, 3504, -157, -3332, -115, 3150, 
396, -2950, -688, 2746, 988, -2526, -1285, 2295, 1590, 
-2050, -1889, 1801, 2179, -1558, -2489, 1308, 2772, -1069, 
-3061, 811, 3344, -575, -3605, 337, 3847, -110, -4095, 
-122, 4317, 325, -4521, -535, 4705, 710, -4881, -888, 
5034, 1047, -5165, -1186, 5263, 1300, -5363, -1409, 5432, 
1499, -5468, -1549, 5483, 1601, -5488, -1614, 5479, 1616, 
-5434, -1605, 5377, 1560, -5296, -1500, 5199, 1427, -5067, 
-1325, 4947, 1193, -4796, -1070, 4624, 911, -4461, -752, 
4267, 564, -4078, -368, 3869, 168, -3649, 59, 3436, 
-276, -3224, 510, 3004, -750, -2780, 986, 2549, -1214, 
-2344, 1454, 2125, -1698, -1905, 1935, 1712, -2160, -1510, 
2378, 1327, -2589, -1156, 2791, 999, -2971, -853, 3142, 
711, -3314, -593, 3455, 477, -3576, -387, 3693, 310, 
-3772, -239, 3855, 189, -3896, -155, 3926, 140, -3930, 
-150, 3924, 154, -3897, -181, 3835, 236, -3767, -284, 
3670, 343, -3558, -427, 3419, 523, -3281, -618, 3107, 
724, -2938, -846, 2743, 969, -2533, -1090, 2316, 1226, 
-2090, -1358, 1854, 1486, -1602, -1631, 1366, 1770, -1110, 
-1908, 859, 2038, -603, -2174, 354, 2305, -113, -2423, 
-133, 2543, 375, -2656, -599, 2748, 808, -2841, -1017, 
2934, 1214, -3007, -1390, 3078, 1557, -3128, -1704, 3179, 
1852, -3224, -1955, 3247, 2053, -3273, -2141, 3278, 2212, 
-3278, -2248, 3266, 2268, -3235, -2289, 3209, 2272, -3165, 
-2244, 3129, 2198, -3068, -2130, 3020, 2058, -2946, -1970, 
2886, 1864, -2813, -1746, 2732, 1607, -2642, -1458, 2559, 
1309, -2475, -1162, 2384, 1001, -2303, -832, 2204, 662, 
-2123, -489, 2036, 320, -1950, -154, 1875, -21, -1792, 
174, 1711, -324, -1638, 472, 1584, -620, -1505, 747, 
1461, -853, -1394, 967, 1341, -1057, -1308, 1133, 1260, 
-1192, -1225, 1239, 1199, -1273, -1160, 1296, 1135, -1294, 
-1126, 1275, 1102, -1247, -1093, 1198, 1065, -1134, -1056, 
1050, 1046, -961, -1050, 851, 1041, -739, -1016, 609, 
1018, -461, -1009, 319, 997, -165, -979, 8, 955, 
164, -941, -322, 915, 498, -879, -660, 853, 835, 
-808, -1002, 766, 1164, -725, -1320, 671, 1453, -607, 
-1588, 555, 1724, -471, -1838, 397, 1931, -317, -2021, 
245, 2088, -144, -2136, 56, 2182, 37, -2199, -146, 
2188, 246, -2172, -358, 2136, 481, -2078, -594, 1990, 
705, -1895, -824, 1777, 947, -1638, -1067, 1480, 1181, 
-1317, -1296, 1130, 1415, -919, -1514, 710, 1627, -477, 
-1729, 235, 1839, 20, -1936, -283, 2013, 547, -2104, 
-808, 2173, 1091, -2244, -1373, 2310, 1640, -2372, -1908, 
2415, 2185, -2459, -2454, 2487, 2697, -2503, -2952, 2513, 
3181, -2517, -3395, 2504, 3614, -2486, -3804, 2468, 3979, 
-2433, -4126, 2379, 4263, -2332, -4379, 2275, 4466, -2196, 
-4535, 2116, 4571, -2028, -4604, 1948, 4599, -1839, -4560, 
1735, 4518, -1622, -4437, 1501, 4336, -1394, -4210, 1266, 
4067, -1122, -3888, 1003, 3696, -865, -3496, 726, 3265, 
-586, -3012, 450, 2757, -311, -2471, 155, 2178, -29, 
-1867, -109, 1554, 256, -1230, -394, 908, 524, -577, 
-644, 239, 765, 100, -885, -436, 1005, 770, -1120, 
-1093, 1230, 1416, -1334, -1734, 1426, 2045, -1516, -2351, 
1589, 2625, -1672, -2894, 1742, 3161, -1800, -3398, 1861, 
3625, -1909, -3828, 1947, 4024, -1967, -4195, 2004, 4349, 
-2008, -4475, 2023, 4598, -2019, -4696, 2027, 4775, -2001, 
-4834, 1980, 4876, -1957, -4907, 1917, 4909, -1864, -4909, 
1821, 4877, -1761, -4852, 1688, 4798, -1622, -4745, 1530, 
4666, -1443, -4594, 1358, 4514, -1246, -4416, 1136, 4316, 
-1025, -4220, 914, 4117, -779, -4021, 657, 3913, -529, 
-3819, 389, 3720, -239, -3630, 87, 3548, 52, -3461, 
-202, 3379, 355, -3318, -515, 3264, 681, -3216, -836, 
3181, 991, -3154, -1143, 3136, 1302, -3125, -1455, 3126, 
1602, -3138, -1745, 3163, 1889, -3187, -2035, 3228, 2162, 
-3280, -2294, 3347, 2408, -3404, -2515, 3481, 2630, -3557, 
-2722, 3625, 2812, -3716, -2884, 3799, 2951, -3882, -2998, 
3953, 3046, -4042, -3071, 4120, 3086, -4194, -3096, 4258, 
3084, -4321, -3061, 4370, 3032, -4406, -2976, 4429, 2913, 
-4450, -2844, 4467, 2749, -4452, -2654, 4430, 2536, -4397, 
-2413, 4344, 2271, -4293, -2129, 4210, 1965, -4101, -1813, 
3991, 1630, -3864, -1446, 3723, 1258, -3550, -1055, 3385, 
858, -3181, -654, 2990, 448, -2765, -241, 2539, 42, 
-2293, 164, 2045, -366, -1785, 558, 1516, -741, -1234, 
930, 967, -1099, -674, 1266, 398, -1416, -114, 1568, 
-179, -1693, 462, 1809, -741, -1893, 1012, 1981, -1273, 
-2045, 1528, 2093, -1773, -2121, 2010, 2113, -2227, -2104, 
2437, 2065, -2633, -2018, 2820, 1931, -2979, -1841, 3128, 
1725, -3251, -1590, 3370, 1425, -3458, -1246, 3532, 1050, 
-3594, -847, 3632, 618, -3650, -372, 3642, 118, -3617, 
154, 3592, -439, -3544, 735, 3470, -1029, -3388, 1329, 
3283, -1647, -3174, 1965, 3053, -2281, -2909, 2591, 2776, 
-2901, -2619, 3208, 2446, -3508, -2287, 3807, 2112, -4083, 
-1935, 4348, 1765, -4606, -1585, 4848, 1406, -5063, -1243, 
5269, 1073, -5444, -891, 5619, 743, -5751, -578, 5867, 
438, -5952, -290, 6020, 170, -6065, -46, 6076, -55, 
-6057, 156, 6031, -255, -5967, 317, 5875, -386, -5757, 
436, 5610, -484, -5449, 513, 5257, -524, -5048, 533, 
4816, -540, -4554, 525, 4292, -508, -4001, 472, 3707, 
-434, -3385, 385, 3053, -349, -2722, 293, 2392, -225, 
-2044, 167, 1685, -107, -1334, 41, 987, 19, -645, 
-78, 314, 138, 26, -194, -340, 241, 659, -286, 
-942, 328, 1224, -367, -1497, 381, 1745, -414, -1968, 
412, 2176, -415, -2366, 408, 2530, -396, -2660, 363, 
2771, -314, -2869, 281, 2927, -211, -2974, 159, 2997, 
-76, -2994, 0, 2960, 93, -2906, -199, 2835, 300, 
-2732, -413, 2610, 527, -2473, -641, 2333, 770, -2150, 
-885, 1965, 1016, -1774, -1131, 1577, 1258, -1356, -1378, 
1130, 1498, -903, -1619, 675, 1723, -436, -1824, 211, 
1918, 26, -2004, -254, 2069, 463, -2134, -678, 2182, 
888, -2234, -1077, 2266, 1249, -2275, -1424, 2275, 1575, 
-2262, -1697, 2245, 1812, -2194, -1912, 2145, 2005, -2081, 
-2067, 1999, 2099, -1887, -2129, 1783, 2117, -1660, -2112, 
1514, 2069, -1365, -2007, 1211, 1936, -1031, -1856, 863, 
1748, -671, -1612, 460, 1476, -257, -1330, 49, 1165, 
171, -994, -392, 806, 621, -618, -852, 419, 1072, 
-226, -1308, 28, 1523, 185, -1746, -372, 1964, 579, 
-2188, -768, 2391, 967, -2592, -1137, 2790, 1313, -2968, 
-1474, 3146, 1623, -3318, -1751, 3466, 1877, -3615, -1983, 
3751, 2081, -3863, -2161, 3971, 2217, -4078, -2264, 4155, 
2286, -4231, -2289, 4288, 2272, -4328, -2237, 4358, 2192, 
-4388, -2128, 4393, 2044, -4392, -1947, 4372, 1833, -4352, 
-1703, 4311, 1573, -4268, -1419, 4218, 1250, -4149, -1074, 
4070, 895, -3992, -698, 3905, 510, -3799, -305, 3709, 
113, -3593, 84, 3493, -301, -3379, 495, 3257, -696, 
-3136, 879, 3002, -1073, -2880, 1244, 2757, -1412, -2627, 
1577, 2483, -1733, -2361, 1870, 2232, -1993, -2089, 2107, 
1955, -2213, -1831, 2292, 1709, -2367, -1567, 2420, 1440, 
-2466, -1313, 2482, 1196, -2504, -1059, 2497, 935, -2474, 
-826, 2445, 693, -2392, -582, 2341, 467, -2267, -346, 
2181, 217, -2075, -117, 1981, -4, -1873, 111, 1746, 
-216, -1622, 325, 1482, -435, -1346, 549, 1216, -639, 
-1060, 747, 922, -828, -785, 933, 631, -1012, -493, 
1095, 356, -1178, -219, 1256, 102, -1320, 27, 1373, 
-152, -1437, 262, 1480, -360, -1524, 451, 1555, -551, 
-1569, 622, 1584, -695, -1584, 763, 1579, -820, -1550, 
851, 1520, -887, -1481, 919, 1411, -951, -1351, 964, 
1268, -972, -1158, 972, 1043, -951, -914, 948, 785, 
-937, -623, 919, 462, -893, -274, 861, 74, -833, 
127, 803, -354, -772, 600, 756, -845, -719, 1105, 
695, -1373, -678, 1639, 655, -1926, -633, 2224, 621, 
-2512, -611, 2814, 610, -3117, -608, 3421, 620, -3730, 
-635, 4026, 646, -4331, -667, 4637, 694, -4930, -726, 
5200, 767, -5485, -810, 5743, 856, -5989, -901, 6229, 
949, -6456, -1007, 6659, 1060, -6845, -1124, 7012, 1192, 
-7156, -1252, 7279, 1302, -7381, -1373, 7457, 1424, -7514, 
-1491, 7545, 1538, -7535, -1584, 7515, 1638, -7479, -1675, 
7397, 1718, -7307, -1754, 7170, 1771, -7032, -1791, 6858, 
1805, -6660, -1819, 6445, 1826, -6192, -1819, 5933, 1805, 
-5644, -1782, 5345, 1755, -5043, -1705, 4711, 1677, -4371, 
-1614, 4009, 1564, -3651, -1499, 3275, 1430, -2899, -1356, 
2521, 1280, -2128, -1197, 1750, 1116, -1385, -1033, 1009, 
939, -645, -845, 294, 758, 57, -663, -385, 578, 
703, -470, -992, 386, 1273, -302, -1540, 218, 1771, 
-136, -1999, 53, 2181, 22, -2345, -103, 2502, 159, 
-2607, -228, 2704, 293, -2766, -332, 2798, 385, -2807, 
-431, 2799, 472, -2745, -499, 2684, 527, -2587, -552, 
2480, 565, -2332, -593, 2171, 593, -1990, -602, 1782, 
609, -1564, -629, 1334, 631, -1082, -640, 823, 642, 
-547, -633, 276, 643, 10, -650, -306, 667, 590, 
-684, -890, 692, 1162, -708, -1451, 733, 1728, -765, 
-1990, 796, 2260, -833, -2499, 885, 2721, -927, -2943, 
978, 3141, -1049, -3309, 1111, 3469, -1186, -3606, 1260, 
3704, -1339, -3797, 1413, 3863, -1498, -3901, 1595, 3919, 
-1686, -3902, 1770, 3862, -1867, -3806, 1957, 3713, -2058, 
-3589, 2148, 3449, -2232, -3298, 2311, 3115, -2386, -2902, 
2462, 2674, -2529, -2416, 2591, 2162, -2633, -1873, 2676, 
1577, -2701, -1254, 2713, 939, -2718, -600, 2710, 246, 
-2689, 94, 2658, -453, -2613, 809, 2543, -1163, -2466, 
1527, 2371, -1887, -2265, 2235, 2146, -2576, -2015, 2912, 
1864, -3243, -1686, 3563, 1511, -3856, -1334, 4155, 1122, 
-4426, -925, 4684, 702, -4923, -476, 5145, 240, -5332, 
2, 5524, -252, -5686, 495, 5818, -734, -5936, 989, 
6043, -1227, -6119, 1478, 6172, -1702, -6197, 1931, 6215, 
-2157, -6210, 2373, 6172, -2572, -6133, 2768, 6053, -2943, 
-5977, 3101, 5870, -3236, -5763, 3365, 5634, -3475, -5488, 
3576, 5329, -3641, -5159, 3698, 4981, -3723, -4791, 3731, 
4583, -3727, -4390, 3702, 4183, -3651, -3977, 3571, 3755, 
-3484, -3544, 3374, 3346, -3260, -3127, 3111, 2914, -2957, 
-2715, 2795, 2516, -2601, -2323, 2414, 2135, -2208, -1953, 
1998, 1773, -1782, -1608, 1557, 1451, -1342, -1318, 1123, 
1180, -898, -1057, 686, 949, -480, -836, 263, 746, 
-68, -669, -101, 606, 281, -543, -421, 500, 567, 
-453, -682, 429, 781, -417, -869, 403, 926, -407, 
-966, 419, 981, -436, -970, 474, 938, -506, -887, 
531, 804, -584, -710, 633, 579, -675, -438, 731, 
259, -788, -77, 847, -134, -900, 365, 948, -605, 
-1007, 867, 1071, -1140, -1118, 1421, 1175, -1724, -1208, 
2016, 1261, -2327, -1299, 2639, 1333, -2951, -1347, 3257, 
1381, -3555, -1383, 3870, 1396, -4160, -1397, 4435, 1382, 
-4712, -1366, 4962, 1351, -5205, -1316, 5417, 1266, -5615, 
-1223, 5793, 1170, -5939, -1099, 6082, 1022, -6180, -938, 
6251, 861, -6303, -757, 6326, 652, -6315, -532, 6265, 
409, -6198, -285, 6104, 150, -5973, -16, 5824, -134, 
-5643, 273, 5423, -423, -5197, 585, 4938, -750, -4649, 
908, 4348, -1083, -4033, 1250, 3690, -1410, -3339, 1590, 
2959, -1749, -2587, 1911, 2197, -2087, -1810, 2237, 1398, 
-2401, -1009, 2558, 613, -2705, -202, 2853, -188, -2987, 
562, 3128, -947, -3251, 1309, 3360, -1653, -3463, 1981, 
3567, -2307, -3644, 2603, 3728, -2870, -3784, 3123, 3850, 
-3349, -3888, 3555, 3908, -3743, -3926, 3900, 3935, -4017, 
-3923, 4124, 3880, -4196, -3842, 4249, 3799, -4270, -3724, 
4264, 3631, -4227, -3539, 4181, 3423, -4097, -3296, 3996, 
3157, -3868, -3004, 3736, 2837, -3568, -2652, 3388, 2452, 
-3195, -2247, 2989, 2036, -2773, -1793, 2540, 1569, -2301, 
-1316, 2062, 1062, -1822, -808, 1568, 533, -1323, -258, 
1070, -20, -820, 286, 597, -577, -365, 856, 128, 
-1131, 69, 1419, -271, -1678, 462, 1952, -644, -2222, 
792, 2472, -935, -2733, 1060, 2957, -1184, -3197, 1275, 
3415, -1342, -3615, 1403, 3811, -1441, -3974, 1456, 4131, 
-1461, -4276, 1442, 4407, -1405, -4506, 1363, 4594, -1291, 
-4669, 1226, 4707, -1131, -4741, 1030, 4749, -913, -4720, 
780, 4696, -654, -4643, 505, 4566, -348, -4464, 205, 
4348, -49, -4205, -122, 4054, 279, -3874, -445, 3680, 
601, -3473, -758, 3234, 901, -2997, -1051, 2746, 1201, 
-2465, -1337, 2197, 1465, -1904, -1578, 1593, 1692, -1290, 
-1777, 980, 1875, -667, -1948, 339, 2016, -6, -2064, 
-318, 2113, 631, -2130, -960, 2160, 1280, -2167, -1596, 
2161, 1889, -2141, -2191, 2111, 2481, -2081, -2763, 2038, 
3030, -1984, -3289, 1919, 3531, -1843, -3750, 1768, 3966, 
-1690, -4171, 1613, 4341, -1513, -4512, 1415, 4663, -1327, 
-4795, 1222, 4903, -1117, -4986, 1017, 5065, -927, -5119, 
826, 5175, -728, -5193, 626, 5196, -534, -5193, 439, 
5171, -364, -5121, 280, 5073, -190, -5005, 120, 4926, 
-62, -4832, -4, 4732, 61, -4609, -121, 4489, 169, 
-4367, -213, 4219, 245, -4075, -269, 3935, 302, -3789, 
-319, 3630, 349, -3475, -358, 3327, 369, -3172, -394, 
3025, 396, -2876, -403, 2720, 404, -2577, -404, 2440, 
411, -2309, -405, 2174, 412, -2047, -409, 1942, 401, 
-1829, -414, 1723, 413, -1627, -419, 1541, 423, -1469, 
-429, 1388, 427, -1335, -443, 1274, 442, -1221, -468, 
1173, 467, -1137, -491, 1104, 506, -1074, -515, 1057, 
528, -1038, -551, 1016, 566, -1005, -587, 992, 609, 
-985, -617, 977, 632, -976, -660, 957, 668, -961, 
-674, 943, 685, -933, -687, 930, 684, -909, -691, 
902, 685, -867, -682, 839, 661, -817, -641, 784, 
635, -751, -594, 695, 579, -651, -536, 601, 494, 
-554, -455, 492, 414, -420, -361, 358, 290, -279, 
-245, 211, 178, -127, -115, 56, 42, 29, 31, 
-109, -102, 200, 187, -272, -256, 360, 346, -432, 
-425, 511, 508, -596, -584, 661, 667, -734, -744, 
789, 826, -860, -893, 907, 980, -955, -1044, 987, 
1116, -1016, -1172, 1039, 1247, -1063, -1301, 1073, 1364, 
-1069, -1409, 1052, 1464, -1028, -1512, 1011, 1550, -976, 
-1588, 928, 1616, -860, -1659, 802, 1687, -728, -1699, 
649, 1724, -550, -1753, 448, 1770, -343, -1780, 231, 
1800, -115, -1810, -2, 1822, 135, -1842, -263, 1853, 
398, -1868, -536, 1879, 667, -1904, -809, 1919, 947, 
-1940, -1092, 1960, 1232, -1995, -1367, 2015, 1507, -2053, 
-1641, 2085, 1761, -2124, -1881, 2171, 2004, -2229, -2119, 
2278, 2212, -2338, -2318, 2398, 2409, -2453, -2483, 2526, 
2571, -2581, -2634, 2662, 2701, -2741, -2748, 2804, 2798, 
-2885, -2829, 2957, 2849, -3045, -2879, 3121, 2886, -3199, 
-2892, 3269, 2884, -3347, -2876, 3404, 2849, -3483, -2824, 
3544, 2798, -3602, -2773, 3640, 2724, -3696, -2685, 3738, 
2636, -3755, -2585, 3788, 2536, -3795, -2478, 3808, 2416, 
-3803, -2344, 3788, 2289, -3761, -2222, 3717, 2161, -3680, 
-2104, 3620, 2038, -3554, -1978, 3469, 1911, -3377, -1860, 
3277, 1800, -3176, -1738, 3054, 1686, -2914, -1630, 2786, 
1574, -2635, -1520, 2478, 1472, -2320, -1414, 2140, 1377, 
-1967, -1327, 1787, 1278, -1599, -1229, 1406, 1168, -1219, 
-1117, 1014, 1070, -821, -1016, 616, 953, -426, -899, 
220, 833, -25, -758, -164, 687, 350, -621, -533, 
533, 714, -448, -877, 370, 1050, -276, -1208, 182, 
1358, -63, -1510, -48, 1653, 151, -1775, -271, 1893, 
409, -2008, -532, 2100, 675, -2198, -806, 2295, 949, 
-2361, -1093, 2439, 1244, -2496, -1401, 2534, 1545, -2583, 
-1690, 2627, 1855, -2657, -2001, 2684, 2149, -2693, -2286, 
2703, 2426, -2708, -2557, 2721, 2689, -2723, -2807, 2721, 
2914, -2713, -3007, 2702, 3111, -2704, -3175, 2688, 3237, 
-2678, -3292, 2674, 3334, -2673, -3357, 2660, 3358, -2667, 
-3341, 2655, 3305, -2651, -3259, 2665, 3192, -2668, -3106, 
2674, 3001, -2678, -2866, 2685, 2729, -2708, -2560, 2717, 
2370, -2739, -2173, 2758, 1943, -2774, -1709, 2801, 1446, 
-2814, -1179, 2841, 900, -2860, -589, 2877, 275, -2881, 
54, 2905, -393, -2904, 738, 2905, -1076, -2912, 1439, 
2905, -1808, -2895, 2171, 2885, -2532, -2868, 2906, 2823, 
-3258, -2800, 3626, 2752, -3973, -2695, 4311, 2629, -4648, 
-2557, 4963, 2477, -5277, -2389, 5556, 2294, -5838, -2179, 
6104, 2067, -6327, -1940, 6554, 1800, -6757, -1656, 6917, 
1510, -7083, -1365, 7208, 1204, -7314, -1022, 7388, 855, 
-7432, -675, 7459, 499, -7462, -318, 7450, 139, -7403, 
39, 7329, -215, -7232, 400, 7104, -569, -6971, 749, 
6806, -898, -6636, 1061, 6428, -1217, -6214, 1355, 5986, 
-1489, -5734, 1613, 5480, -1731, -5220, 1830, 4940, -1920, 
-4661, 1993, 4372, -2060, -4079, 2113, 3786, -2146, -3497, 
2166, 3200, -2158, -2918, 2149, 2640, -2125, -2378, 2090, 
2118, -2026, -1866, 1967, 1624, -1878, -1398, 1785, 1200, 
-1675, -1004, 1563, 825, -1429, -668, 1295, 546, -1136, 
-425, 981, 324, -814, -240, 653, 192, -487, -142, 
300, 129, -124, -128, -53, 144, 224, -180, -411, 
244, 582, -315, -741, 403, 909, -492, -1061, 614, 
1216, -734, -1342, 861, 1467, -1016, -1589, 1167, 1703, 
-1326, -1794, 1477, 1869, -1632, -1940, 1809, 1993, -1965, 
-2022, 2128, 2056, -2272, -2060, 2418, 2051, -2559, -2029, 
2686, 2008, -2819, -1957, 2915, 1887, -3015, -1823, 3093, 
1735, -3164, -1625, 3215, 1517, -3253, -1398, 3268, 1277, 
-3276, -1146, 3257, 1000, -3233, -849, 3181, 692, -3109, 
-551, 3029, 391, -2919, -236, 2806, 62, -2672, 85, 
2527, -244, -2362, 386, 2189, -539, -2008, 671, 1805, 
-798, -1598, 931, 1394, -1041, -1171, 1149, 955, -1242, 
-725, 1320, 507, -1391, -274, 1449, 52, -1510, 155, 
1544, -366, -1562, 586, 1566, -781, -1561, 969, 1536, 
-1146, -1512, 1320, 1472, -1480, -1414, 1616, 1349, -1739, 
-1271, 1861, 1184, -1957, -1073, 2042, 962, -2107, -855, 
2144, 736, -2180, -593, 2197, 465, -2193, -321, 2172, 
188, -2132, -33, 2080, -112, -2010, 262, 1944, -421, 
-1840, 555, 1748, -707, -1636, 850, 1510, -988, -1378, 
1126, 1250, -1259, -1121, 1386, 969, -1500, -835, 1614, 
681, -1708, -547, 1804, 396, -1899, -277, 1987, 136, 
-2057, -29, 2109, -86, -2177, 198, 2223, -290, -2250, 
355, 2291, -429, -2311, 471, 2326, -516, -2325, 530, 
2330, -540, -2324, 525, 2307, -492, -2281, 450, 2262, 
-378, -2235, 303, 2203, -197, -2167, 83, 2120, 38, 
-2070, -176, 2035, 326, -1983, -503, 1930, 677, -1881, 
-867, 1830, 1073, -1781, -1266, 1744, 1486, -1698, -1698, 
1648, 1924, -1602, -2144, 1549, 2357, -1506, -2568, 1462, 
2776, -1432, -2992, 1382, 3187, -1353, -3364, 1308, 3543, 
-1274, -3718, 1239, 3875, -1208, -4003, 1163, 4127, -1126, 
-4232, 1101, 4317, -1059, -4370, 1027, 4428, -987, -4443, 
943, 4445, -906, -4432, 857, 4393, -808, -4323, 758, 
4239, -701, -4129, 641, 3998, -583, -3859, 524, 3677, 
-452, -3499, 377, 3285, -303, -3064, 225, 2818, -138, 
-2576, 36, 2296, 51, -2028, -149, 1733, 259, -1423, 
-357, 1127, 465, -814, -575, 503, 689, -173, -809, 
-138, 912, 455, -1027, -765, 1150, 1083, -1258, -1382, 
1385, 1676, -1495, -1951, 1593, 2226, -1710, -2499, 1814, 
2736, -1905, -2969, 1998, 3198, -2093, -3403, 2164, 3592, 
-2247, -3753, 2303, 3898, -2359, -4039, 2424, 4157, -2461, 
-4254, 2497, 4325, -2513, -4391, 2521, 4434, -2538, -4444, 
2523, 4450, -2511, -4454, 2491, 4424, -2447, -4392, 2411, 
4340, -2355, -4272, 2288, 4200, -2209, -4106, 2127, 4012, 
-2050, -3923, 1954, 3812, -1841, -3691, 1733, 3577, -1613, 
-3454, 1499, 3336, -1372, -3220, 1240, 3087, -1121, -2981, 
989, 2862, -845, -2753, 714, 2632, -573, -2545, 437, 
2448, -303, -2357, 171, 2277, -31, -2190, -84, 2135, 
222, -2070, -337, 2022, 454, -1969, -565, 1939, 672, 
-1899, -775, 1890, 879, -1857, -960, 1853, 1052, -1841, 
-1144, 1849, 1209, -1839, -1284, 1850, 1342, -1843, -1413, 
1850, 1469, -1858, -1516, 1856, 1559, -1855, -1600, 1844, 
1646, -1821, -1683, 1812, 1706, -1775, -1739, 1740, 1775, 
-1693, -1809, 1636, 1836, -1573, -1856, 1493, 1875, -1408, 
-1900, 1301, 1940, -1200, -1961, 1070, 1989, -923, -2021, 
776, 2056, -593, -2079, 422, 2116, -230, -2153, 19, 
2181, 191, -2213, -429, 2253, 658, -2295, -905, 2343, 
1163, -2373, -1418, 2419, 1677, -2446, -1944, 2494, 2216, 
-2517, -2482, 2559, 2759, -2579, -3025, 2611, 3292, -2629, 
-3545, 2645, 3798, -2640, -4037, 2639, 4256, -2641, -4474, 
2628, 4665, -2598, -4864, 2571, 5015, -2523, -5167, 2463, 
5306, -2404, -5411, 2332, 5496, -2244, -5544, 2140, 5592, 
-2023, -5598, 1906, 5589, -1759, -5545, 1617, 5491, -1452, 
-5403, 1278, 5287, -1084, -5148, 884, 4985, -670, -4795, 
454, 4583, -225, -4339, -8, 4096, 262, -3818, -497, 
3513, 763, -3217, -1019, 2883, 1281, -2551, -1552, 2194, 
1817, -1828, -2083, 1463, 2340, -1091, -2584, 715, 2845, 
-330, -3081, -52, 3307, 422, -3529, -803, 3743, 1155, 
-3943, -1508, 4121, 1861, -4291, -2186, 4440, 2507, -4566, 
-2807, 4673, 3090, -4770, -3351, 4836, 3588, -4880, -3803, 
4895, 4004, -4899, -4170, 4879, 4311, -4827, -4430, 4749, 
4520, -4654, -4576, 4528, 4628, -4398, -4641, 4224, 4617, 
-4033, -4585, 3829, 4514, -3591, -4413, 3346, 4301, -3081, 
-4173, 2793, 4016, -2501, -3835, 2184, 3637, -1861, -3422, 
1541, 3201, -1188, -2947, 852, 2702, -499, -2443, 142, 
2159, 202, -1894, -553, 1616, 912, -1322, -1260, 1038, 
1580, -771, -1911, 487, 2225, -220, -2523, -37, 2813, 
291, -3078, -527, 3336, 762, -3567, -975, 3784, 1166, 
-3971, -1350, 4144, 1521, -4289, -1662, 4407, 1785, -4509, 
-1886, 4580, 1976, -4624, -2040, 4648, 2071, -4639, -2105, 
4615, 2104, -4561, -2086, 4479, 2043, -4383, -1984, 4250, 
1909, -4112, -1816, 3941, 1700, -3767, -1580, 3563, 1437, 
-3355, -1294, 3133, 1135, -2877, -964, 2632, 774, -2370, 
-595, 2115, 395, -1841, -212, 1558, 7, -1290, 187, 
1005, -377, -726, 568, 468, -748, -195, 918, -62, 
-1097, 305, 1246, -546, -1394, 769, 1545, -992, -1671, 
1181, 1776, -1378, -1879, 1534, 1944, -1690, -2020, 1825, 
2070, -1936, -2095, 2041, 2117, -2111, -2113, 2172, 2092, 
-2209, -2061, 2239, 2003, -2237, -1946, 2215, 1867, -2179, 
-1765, 2133, 1661, -2081, -1550, 1996, 1422, -1909, -1277, 
1789, 1122, -1676, -965, 1545, 817, -1422, -638, 1270, 
474, -1126, -307, 968, 132, -806, 38, 648, -189, 
-481, 351, 324, -507, -159, 666, 4, -794, 145, 
932, -284, -1045, 426, 1155, -549, -1245, 670, 1331, 
-782, -1389, 885, 1445, -989, -1491, 1054, 1509, -1131, 
-1500, 1187, 1500, -1232, -1470, 1264, 1425, -1282, -1365, 
1272, 1284, -1272, -1188, 1263, 1088, -1225, -969, 1187, 
833, -1144, -690, 1082, 528, -1010, -365, 934, 202, 
-855, -15, 765, -168, -673, 365, 572, -556, -483, 
748, 376, -943, -274, 1145, 174, -1327, -89, 1521, 
-17, -1698, 109, 1875, -183, -2035, 261, 2192, -341, 
-2347, 403, 2485, -465, -2607, 519, 2723, -552, -2818, 
582, 2891, -601, -2958, 602, 3019, -601, -3057, 585, 
3061, -559, -3072, 517, 3057, -475, -3029, 406, 2982, 
-324, -2924, 254, 2843, -159, -2764, 47, 2659, 61, 
-2548, -183, 2423, 322, -2275, -457, 2128, 600, -1980, 
-761, 1830, 904, -1656, -1066, 1500, 1242, -1316, -1406, 
1157, 1577, -979, -1742, 813, 1917, -649, -2087, 488, 
2253, -325, -2418, 181, 2589, -50, -2741, -86, 2910, 
200, -3051, -314, 3207, 406, -3347, -492, 3483, 555, 
-3610, -595, 3729, 634, -3855, -652, 3957, 662, -4061, 
-636, 4159, 610, -4246, -564, 4324, 511, -4388, -428, 
4448, 340, -4517, -232, 4570, 105, -4613, 16, 4641, 
-169, -4683, 309, 4710, -483, -4722, 656, 4752, -829, 
-4760, 1014, 4756, -1197, -4761, 1387, 4761, -1571, -4763, 
1765, 4745, -1950, -4745, 2135, 4722, -2314, -4716, 2478, 
4692, -2648, -4668, 2794, 4651, -2941, -4625, 3070, 4589, 
-3178, -4567, 3270, 4526, -3361, -4493, 3418, 4452, -3467, 
-4407, 3497, 4372, -3500, -4312, 3481, 4270, -3456, -4213, 
3388, 4146, -3323, -4078, 3223, 4013, -3109, -3936, 2974, 
3860, -2819, -3779, 2632, 3672, -2441, -3583, 2236, 3475, 
-2004, -3355, 1766, 3236, -1508, -3109, 1248, 2972, -968, 
-2826, 678, 2674, -379, -2507, 79, 2341, 231, -2155, 
-527, 1967, 845, -1765, -1142, 1567, 1449, -1359, -1754, 
1133, 2047, -921, -2322, 692, 2605, -446, -2867, 206, 
3108, 35, -3347, -285, 3569, 533, -3768, -799, 3950, 
1056, -4111, -1308, 4242, 1560, -4351, -1824, 4455, 2066, 
-4518, -2329, 4576, 2571, -4598, -2802, 4600, 3052, -4573, 
-3278, 4521, 3498, -4459, -3708, 4356, 3904, -4249, -4101, 
4116, 4277, -3944, -4451, 3783, 4611, -3584, -4762, 3369, 
4894, -3155, -5018, 2907, 5126, -2657, -5212, 2405, 5282, 
-2127, -5353, 1860, 5391, -1582, -5429, 1296, 5452, -1014, 
-5458, 744, 5441, -467, -5426, 195, 5384, 67, -5327, 
-328, 5274, 568, -5205, -803, 5131, 1020, -5039, -1223, 
4929, 1400, -4825, -1578, 4719, 1714, -4597, -1849, 4475, 
1954, -4350, -2032, 4214, 2097, -4088, -2129, 3956, 2139, 
-3814, -2141, 3689, 2099, -3571, -2044, 3447, 1965, -3329, 
-1881, 3212, 1754, -3109, -1614, 3017, 1460, -2916, -1292, 
2839, 1098, -2766, -883, 2701, 670, -2663, -447, 2623, 
193, -2591, 45, 2583, -295, -2563, 558, 2578, -811, 
-2598, 1081, 2626, -1328, -2663, 1582, 2730, -1829, -2782, 
2062, 2865, -2301, -2954, 2519, 3051, -2713, -3155, 2900, 
3260, -3070, -3383, 3215, 3495, -3360, -3634, 3454, 3774, 
-3545, -3915, 3623, 4052, -3659, -4195, 3682, 4344, -3670, 
-4478, 3635, 4619, -3576, -4768, 3502, 4904, -3387, -5040, 
3255, 5171, -3100, -5285, 2919, 5399, -2734, -5513, 2501, 
5611, -2277, -5685, 2015, 5773, -1740, -5831, 1462, 5895, 
-1163, -5933, 852, 5966, -522, -5977, 202, 5984, 125, 
-5975, -461, 5955, 797, -5920, -1128, 5861, 1452, -5808, 
-1767, 5727, 2086, -5626, -2387, 5532, 2679, -5412, -2955, 
5270, 3209, -5136, -3443, 4984, 3662, -4815, -3860, 4631, 
4051, -4447, -4200, 4256, 4326, -4056, -4427, 3848, 4509, 
-3627, -4566, 3398, 4587, -3179, -4585, 2936, 4543, -2717, 
-4497, 2469, 4407, -2240, -4304, 1994, 4170, -1764, -4009, 
1538, 3814, -1309, -3622, 1078, 3396, -855, -3149, 628, 
2877, -422, -2604, 221, 2313, -28, -2011, -163, 1706, 
327, -1378, -499, 1049, 665, -726, -805, 394, 933, 
-58, -1062, -269, 1167, 598, -1256, -902, 1339, 1206, 
-1411, -1511, 1463, 1791, -1496, -2061, 1531, 2306, -1540, 
-2544, 1534, 2756, -1530, -2953, 1502, 3113, -1461, -3275, 
1406, 3393, -1341, -3497, 1264, 3585, -1166, -3629, 1066, 
3669, -946, -3662, 828, 3648, -697, -3617, 563, 3543, 
-411, -3469, 258, 3362, -102, -3231, -74, 3076, 232, 
-2925, -407, 2732, 582, -2552, -769, 2330, 945, -2115, 
-1112, 1895, 1288, -1651, -1462, 1422, 1641, -1177, -1795, 
924, 1959, -676, -2110, 422, 2269, -189, -2406, -44, 
2535, 285, -2651, -510, 2766, 724, -2861, -913, 2943, 
1103, -3014, -1279, 3063, 1443, -3122, -1597, 3139, 1721, 
-3161, -1831, 3160, 1926, -3153, -2011, 3109, 2060, -3069, 
-2111, 3000, 2133, -2922, -2138, 2832, 2129, -2722, -2091, 
2594, 2052, -2458, -1991, 2309, 1919, -2141, -1824, 1963, 
1722, -1769, -1616, 1564, 1504, -1346, -1364, 1114, 1242, 
-881, -1099, 638, 951, -402, -799, 138, 653, 119, 
-497, -369, 361, 639, -210, -907, 70, 1163, 63, 
-1424, -195, 1678, 311, -1935, -422, 2179, 526, -2414, 
-626, 2642, 692, -2853, -764, 3059, 820, -3244, -876, 
3424, 911, -3598, -922, 3739, 930, -3870, -935, 3979, 
913, -4081, -892, 4149, 852, -4215, -790, 4254, 738, 
-4261, -666, 4266, 601, -4241, -517, 4187, 429, -4114, 
-346, 4037, 242, -3922, -144, 3790, 50, -3658, 50, 
3481, -135, -3306, 236, 3097, -322, -2887, 409, 2649, 
-482, -2403, 561, 2160, -627, -1893, 680, 1603, -711, 
-1317, 758, 1033, -773, -726, 778, 425, -784, -117, 
767, -193, -748, 501, 724, -804, -668, 1096, 611, 
-1395, -539, 1693, 467, -1965, -387, 2236, 294, -2508, 
-184, 2751, 68, -3000, 33, 3211, -154, -3429, 273, 
3628, -391, -3803, 516, 3964, -643, -4106, 757, 4223, 
-868, -4338, 971, 4418, -1076, -4495, 1157, 4546, -1241, 
-4575, 1304, 4585, -1366, -4589, 1389, 4570, -1425, -4537, 
1431, 4482, -1415, -4415, 1377, 4345, -1331, -4240, 1274, 
4151, -1168, -4033, 1075, 3900, -943, -3782, 778, 3643, 
-619, -3491, 429, 3343, -216, -3202, -9, 3037, 252, 
-2892, -517, 2745, 797, -2593, -1097, 2450, 1397, -2305, 
-1718, 2170, 2044, -2033, -2376, 1917, 2711, -1813, -3063, 
1714, 3409, -1617, -3749, 1534, 4095, -1469, -4448, 1400, 
4783, -1365, -5110, 1327, 5419, -1298, -5732, 1301, 6023, 
-1298, -6306, 1317, 6572, -1346, -6813, 1375, 7035, -1435, 
-7231, 1482, 7412, -1558, -7573, 1639, 7700, -1717, -7802, 
1818, 7884, -1909, -7931, 2018, 7962, -2132, -7961, 2238, 
7934, -2349, -7877, 2462, 7793, -2577, -7691, 2700, 7544, 
-2809, -7402, 2918, 7227, -3022, -7014, 3115, 6807, -3209, 
-6559, 3295, 6316, -3372, -6036, 3438, 5765, -3486, -5463, 
3534, 5163, -3585, -4848, 3595, 4534, -3626, -4211, 3629, 
3891, -3622, -3565, 3593, 3254, -3565, -2935, 3516, 2627, 
-3468, -2327, 3399, 2035, -3322, -1759, 3244, 1491, -3146, 
-1230, 3038, 991, -2931, -770, 2798, 557, -2678, -358, 
2544, 193, -2403, -47, 2257, -95, -2112, 220, 1952, 
-307, -1812, 395, 1657, -459, -1500, 495, 1335, -532, 
-1198, 542, 1038, -540, -893, 524, 755, -500, -613, 
454, 482, -408, -343, 351, 223, -295, -120, 228, 
12, -154, 90, 83, -188, -14, 286, -42, -367, 
107, 439, -180, -504, 227, 557, -268, -617, 306, 
654, -336, -693, 341, 732, -348, -753, 340, 786, 
-311, -807, 267, 820, -207, -838, 136, 851, -41, 
-852, -52, 867, 183, -864, -312, 882, 460, -886, 
-634, 899, 804, -906, -1002, 913, 1214, -932, -1431, 
947, 1645, -961, -1880, 993, 2123, -1010, -2371, 1044, 
2612, -1084, -2863, 1106, 3117, -1157, -3359, 1196, 3598, 
-1242, -3830, 1287, 4074, -1335, -4283, 1370, 4493, -1420, 
-4705, 1485, 4883, -1530, -5048, 1581, 5206, -1622, -5344, 
1662, 5451, -1712, -5559, 1735, 5633, -1769, -5686, 1804, 
5710, -1829, -5723, 1832, 5707, -1835, -5675, 1844, 5609, 
-1836, -5535, 1812, 5431, -1783, -5312, 1731, 5154, -1690, 
-4990, 1622, 4818, -1548, -4612, 1473, 4398, -1377, -4170, 
1264, 3912, -1146, -3666, 1026, 3401, -877, -3115, 736, 
2831, -570, -2558, 411, 2265, -232, -1967, 68, 1690, 
120, -1405, -311, 1125, 506, -851, -694, 579, 887, 
-321, -1084, 85, 1271, 155, -1464, -361, 1642, 559, 
-1824, -756, 1988, 909, -2144, -1061, 2292, 1184, -2431, 
-1297, 2553, 1388, -2670, -1448, 2754, 1489, -2827, -1512, 
2888, 1518, -2932, -1509, 2952, 1474, -2955, -1415, 2929, 
1342, -2895, -1258, 2834, 1146, -2734, -1023, 2642, 892, 
-2504, -738, 2357, 572, -2194, -411, 2005, 227, -1794, 
-38, 1561, -148, -1328, 336, 1071, -543, -796, 746, 
502, -931, -196, 1133, -113, -1313, 424, 1503, -739, 
-1687, 1082, 1854, -1397, -2022, 1739, 2171, -2069, -2317, 
2398, 2441, -2705, -2553, 3023, 2671, -3328, -2753, 3624, 
2839, -3900, -2900, 4169, 2954, -4409, -2987, 4637, 3016, 
-4846, -3021, 5024, 3014, -5180, -3001, 5324, 2969, -5434, 
-2930, 5513, 2876, -5566, -2811, 5600, 2746, -5600, -2680, 
5582, 2590, -5524, -2511, 5449, 2406, -5326, -2325, 5196, 
2213, -5031, -2128, 4841, 2014, -4632, -1926, 4393, 1836, 
-4139, -1738, 3850, 1648, -3558, -1565, 3241, 1491, -2920, 
-1420, 2575, 1350, -2226, -1294, 1864, 1249, -1494, -1195, 
1115, 1166, -738, -1150, 361, 1131, 18, -1126, -376, 
1118, 749, -1127, -1112, 1133, 1453, -1156, -1786, 1190, 
2102, -1219, -2403, 1250, 2689, -1291, -2971, 1349, 3213, 
-1393, -3442, 1433, 3637, -1474, -3832, 1519, 3980, -1563, 
-4122, 1605, 4218, -1643, -4305, 1682, 4366, -1707, -4398, 
1728, 4408, -1727, -4388, 1728, 4349, -1727, -4281, 1707, 
4204, -1678, -4082, 1630, 3970, -1593, -3818, 1530, 3655, 
-1455, -3475, 1356, 3285, -1255, -3088, 1143, 2876, -1030, 
-2647, 895, 2418, -750, -2179, 592, 1937, -432, -1696, 
255, 1444, -72, -1211, -117, 957, 306, -726, -502, 
497, 716, -278, -916, 65, 1124, 151, -1341, -344, 
1536, 518, -1753, -691, 1947, 859, -2137, -1001, 2339, 
1133, -2522, -1252, 2687, 1347, -2857, -1435, 3020, 1504, 
-3151, -1562, 3296, 1604, -3407, -1640, 3519, 1657, -3606, 
-1662, 3685, 1658, -3748, -1640, 3796, 1622, -3822, -1594, 
3841, 1549, -3829, -1505, 3828, 1453, -3799, -1382, 3753, 
1320, -3704, -1266, 3626, 1195, -3547, -1138, 3455, 1068, 
-3365, -1008, 3259, 943, -3145, -890, 3015, 844, -2887, 
-801, 2764, 749, -2618, -730, 2493, 693, -2362, -684, 
2224, 667, -2101, -671, 1977, 661, -1846, -683, 1750, 
699, -1639, -723, 1539, 756, -1469, -809, 1390, 847, 
-1334, -908, 1287, 951, -1247, -1014, 1237, 1080, -1227, 
-1152, 1227, 1216, -1251, -1290, 1293, 1349, -1354, -1419, 
1420, 1473, -1509, -1540, 1605, 1586, -1724, -1634, 1848, 
1683, -1993, -1709, 2137, 1739, -2295, -1746, 2463, 1764, 
-2637, -1748, 2825, 1743, -3024, -1717, 3215, 1669, -3417, 
-1623, 3618, 1562, -3821, -1482, 4018, 1409, -4220, -1308, 
4405, 1188, -4604, -1072, 4785, 928, -4964, -791, 5142, 
644, -5292, -472, 5440, 299, -5592, -125, 5708, -52, 
-5828, 243, 5934, -452, -6008, 639, 6090, -837, -6146, 
1040, 6195, -1250, -6220, 1450, 6226, -1656, -6236, 1846, 
6219, -2044, -6178, 2229, 6144, -2394, -6084, 2578, 6017, 
-2733, -5933, 2896, 5845, -3028, -5744, 3160, 5632, -3291, 
-5514, 3388, 5389, -3495, -5252, 3569, 5124, -3653, -4977, 
3699, 4841, -3745, -4693, 3784, 4546, -3805, -4416, 3803, 
4262, -3797, -4129, 3781, 3991, -3751, -3871, 3714, 3746, 
-3661, -3627, 3603, 3510, -3532, -3396, 3447, 3306, -3372, 
-3211, 3276, 3139, -3176, -3059, 3080, 2990, -2981, -2939, 
2870, 2879, -2768, -2838, 2660, 2807, -2547, -2783, 2456, 
2764, -2341, -2749, 2238, 2742, -2150, -2729, 2052, 2724, 
-1951, -2719, 1869, 2727, -1796, -2732, 1716, 2734, -1648, 
-2735, 1573, 2730, -1511, -2721, 1465, 2710, -1417, -2694, 
1375, 2668, -1329, -2643, 1286, 2593, -1252, -2556, 1226, 
2497, -1201, -2429, 1176, 2355, -1152, -2256, 1127, 2161, 
-1106, -2055, 1079, 1925, -1040, -1790, 1015, 1634, -988, 
-1476, 949, 1297, -907, -1113, 852, 922, -802, -712, 
723, 495, -655, -275, 578, 43, -499, 189, 404, 
-430, -291, 677, 185, -928, -62, 1182, -79, -1436, 
219, 1686, -361, -1928, 520, 2174, -690, -2414, 862, 
2655, -1035, -2887, 1215, 3098, -1405, -3306, 1582, 3504, 
-1780, -3683, 1976, 3852, -2173, -3998, 2367, 4127, -2555, 
-4248, 2725, 4360, -2909, -4427, 3086, 4497, -3253, -4533, 
3408, 4564, -3543, -4569, 3680, 4555, -3802, -4517, 3900, 
4451, -3983, -4387, 4061, 4277, -4117, -4176, 4146, 4043, 
-4157, -3890, 4159, 3727, -4126, -3540, 4076, 3344, -4007, 
-3131, 3914, 2912, -3813, -2688, 3675, 2444, -3526, -2187, 
3355, 1938, -3155, -1687, 2945, 1422, -2725, -1156, 2472, 
885, -2210, -631, 1934, 372, -1651, -120, 1347, -131, 
-1034, 383, 714, -615, -401, 837, 69, -1055, 269, 
1251, -588, -1431, 915, 1617, -1247, -1770, 1558, 1923, 
-1874, -2053, 2161, 2165, -2457, -2264, 2727, 2343, -2990, 
-2414, 3221, 2451, -3439, -2494, 3632, 2506, -3814, -2501, 
3972, 2479, -4101, -2458, 4194, 2418, -4275, -2352, 4316, 
2287, -4340, -2205, 4318, 2106, -4279, -1996, 4217, 1879, 
-4120, -1767, 3993, 1645, -3826, -1498, 3655, 1363, -3439, 
-1223, 3212, 1089, -2949, -944, 2670, 789, -2352, -639, 
2037, 494, -1686, -352, 1319, 225, -950, -93, 552, 
-38, -146, 167, -266, -284, 690, 408, -1118, -510, 
1539, 604, -1979, -700, 2402, 787, -2838, -859, 3257, 
930, -3670, -1003, 4078, 1045, -4463, -1099, 4840, 1141, 
-5221, -1178, 5570, 1210, -5902, -1244, 6215, 1266, -6509, 
-1282, 6779, 1292, -7022, -1317, 7262, 1327, -7456, -1326, 
7643, 1331, -7797, -1345, 7926, 1363, -8017, -1361, 8106, 
1385, -8146, -1398, 8181, 1418, -8182, -1437, 8168, 1459, 
-8128, -1479, 8054, 1522, -7968, -1549, 7870, 1598, -7742, 
-1636, 7598, 1689, -7435, -1743, 7256, 1803, -7062, -1873, 
6859, 1936, -6644, -2000, 6419, 2074, -6189, -2145, 5949, 
2224, -5687, -2312, 5434, 2383, -5189, -2464, 4938, 2556, 
-4675, -2624, 4413, 2698, -4171, -2771, 3907, 2835, -3672, 
-2904, 3430, 2951, -3198, -3012, 2961, 3056, -2742, -3087, 
2536, 3113, -2328, -3126, 2133, 3134, -1965, -3124, 1793, 
3096, -1624, -3071, 1482, 3028, -1339, -2974, 1224, 2912, 
-1103, -2824, 995, 2735, -919, -2625, 832, 2505, -765, 
-2375, 710, 2232, -668, -2068, 636, 1896, -604, -1723, 
589, 1531, -585, -1343, 590, 1135, -611, -918, 634, 
690, -651, -467, 686, 239, -738, -6, 788, -234, 
-844, 475, 908, -709, -966, 943, 1041, -1172, -1129, 
1399, 1205, -1630, -1288, 1844, 1382, -2058, -1477, 2251, 
1568, -2449, -1659, 2621, 1769, -2782, -1870, 2938, 1973, 
-3087, -2075, 3211, 2183, -3316, -2275, 3413, 2379, -3501, 
-2495, 3564, 2588, -3608, -2694, 3629, 2802, -3634, -2909, 
3638, 3003, -3613, -3107, 3574, 3203, -3504, -3290, 3444, 
3383, -3345, -3466, 3235, 3547, -3122, -3637, 2986, 3697, 
-2843, -3768, 2676, 3847, -2514, -3902, 2323, 3957, -2127, 
-3999, 1939, 4047, -1727, -4072, 1513, 4098, -1297, -4115, 
1073, 4135, -835, -4135, 609, 4143, -393, -4132, 160, 
4116, 67, -4088, -287, 4051, 517, -4012, -726, 3956, 
937, -3897, -1142, 3833, 1336, -3756, -1533, 3678, 1714, 
-3582, -1871, 3502, 2045, -3397, -2194, 3283, 2342, -3176, 
-2473, 3070, 2593, -2950, -2698, 2832, 2794, -2710, -2883, 
2586, 2964, -2466, -3040, 2337, 3086, -2204, -3144, 2090, 
3183, -1963, -3207, 1848, 3218, -1736, -3239, 1633, 3232, 
-1528, -3229, 1434, 3216, -1340, -3193, 1267, 3171, -1195, 
-3142, 1127, 3100, -1084, -3068, 1034, 3023, -997, -2969, 
981, 2910, -969, -2858, 969, 2807, -968, -2738, 997, 
2675, -1028, -2619, 1078, 2543, -1134, -2479, 1201, 2414, 
-1274, -2348, 1362, 2286, -1450, -2203, 1552, 2148, -1657, 
-2067, 1773, 1993, -1893, -1925, 2033, 1854, -2156, -1782, 
2293, 1697, -2439, -1626, 2579, 1539, -2713, -1453, 2851, 
1381, -2976, -1289, 3109, 1197, -3240, -1102, 3369, 1019, 
-3472, -912, 3584, 816, -3679, -705, 3770, 597, -3862, 
-477, 3935, 352, -3992, -235, 4039, 119, -4068, 15, 
4089, -141, -4107, 279, 4088, -423, -4077, 559, 4045, 
-706, -4007, 859, 3941, -995, -3873, 1144, 3788, -1294, 
-3705, 1446, 3592, -1582, -3482, 1734, 3350, -1884, -3221, 
2020, 3074, -2159, -2926, 2289, 2771, -2418, -2600, 2529, 
2436, -2654, -2272, 2747, 2096, -2855, -1936, 2946, 1757, 
-3021, -1602, 3093, 1440, -3158, -1277, 3212, 1112, -3238, 
-973, 3262, 838, -3290, -702, 3279, 573, -3266, -466, 
3247, 363, -3218, -273, 3169, 200, -3099, -120, 3021, 
69, -2943, -26, 2834, -3, -2721, 14, 2603, -16, 
-2463, 20, 2331, -6, -2171, -22, 2014, 66, -1853, 
-118, 1673, 169, -1494, -238, 1319, 318, -1133, -399, 
949, 491, -760, -577, 568, 673, -372, -757, 189, 
862, -10, -960, -162, 1055, 344, -1144, -500, 1235, 
660, -1306, -819, 1380, 959, -1451, -1079, 1523, 1204, 
-1567, -1315, 1615, 1409, -1655, -1483, 1677, 1558, -1684, 
-1604, 1681, 1646, -1661, -1676, 1645, 1676, -1601, -1670, 
1558, 1667, -1485, -1637, 1420, 1579, -1326, -1528, 1234, 
1452, -1130, -1379, 1001, 1281, -874, -1184, 751, 1066, 
-600, -954, 460, 821, -305, -688, 145, 536, 16, 
-399, -167, 244, 330, -95, -485, -60, 642, 198, 
-807, -346, 954, 493, -1092, -641, 1223, 783, -1345, 
-899, 1463, 1034, -1582, -1147, 1666, 1259, -1759, -1343, 
1817, 1436, -1876, -1509, 1920, 1565, -1936, -1626, 1957, 
1667, -1950, -1682, 1932, 1690, -1900, -1693, 1857, 1675, 
-1779, -1645, 1709, 1608, -1616, -1557, 1511, 1490, -1390, 
-1405, 1266, 1313, -1127, -1223, 965, 1105, -806, -995, 
648, 865, -474, -740, 287, 587, -98, -456, -86, 
300, 264, -162, -450, 10, 651, 140, -833, -293, 
1019, 445, -1195, -593, 1354, 729, -1536, -861, 1681, 
988, -1828, -1098, 1983, 1205, -2104, -1309, 2221, 1410, 
-2339, -1489, 2433, 1544, -2523, -1607, 2594, 1648, -2665, 
-1676, 2718, 1687, -2755, -1689, 2776, 1670, -2791, -1648, 
2810, 1607, -2809, -1554, 2787, 1481, -2773, -1408, 2748, 
1320, -2718, -1213, 2680, 1099, -2634, -973, 2596, 844, 
-2538, -693, 2497, 542, -2436, -381, 2390, 224, -2352, 
-53, 2313, -113, -2267, 283, 2241, -473, -2202, 648, 
2179, -820, -2180, 990, 2163, -1155, -2167, 1336, 2177, 
-1490, -2208, 1653, 2230, -1805, -2279, 1945, 2323, -2070, 
-2379, 2206, 2445, -2323, -2531, 2424, 2618, -2534, -2702, 
2611, 2800, -2701, -2905, 2767, 3014, -2819, -3129, 2866, 
3234, -2892, -3348, 2919, 3462, -2930, -3580, 2936, 3690, 
-2931, -3791, 2914, 3896, -2900, -3993, 2865, 4075, -2825, 
-4151, 2789, 4208, -2748, -4260, 2680, 4292, -2635, -4313, 
2573, 4316, -2504, -4300, 2445, 4253, -2383, -4211, 2314, 
4134, -2254, -4035, 2178, 3929, -2132, -3785, 2076, 3639, 
-2009, -3459, 1970, 3249, -1919, -3024, 1883, 2787, -1846, 
-2528, 1801, 2251, -1786, -1938, 1764, 1623, -1746, -1294, 
1749, 952, -1738, -593, 1741, 214, -1753, 161, 1756, 
-544, -1776, 946, 1794, -1348, -1828, 1749, 1847, -2154, 
-1872, 2547, 1917, -2944, -1936, 3340, 1972, -3722, -2007, 
4102, 2027, -4456, -2060, 4815, 2081, -5152, -2095, 5474, 
2102, -5764, -2118, 6055, 2123, -6307, -2107, 6558, 2087, 
-6775, -2066, 6967, 2046, -7128, -2004, 7269, 1958, -7401, 
-1896, 7491, 1819, -7556, -1735, 7606, 1645, -7620, -1541, 
7606, 1429, -7572, -1297, 7526, 1157, -7450, -1022, 7357, 
853, -7243, -690, 7094, 523, -6945, -338, 6781, 157, 
-6602, 45, 6402, -244, -6190, 444, 5985, -651, -5764, 
855, 5535, -1071, -5292, 1273, 5068, -1492, -4831, 1694, 
4603, -1895, -4371, 2107, 4151, -2303, -3929, 2483, 3718, 
-2659, -3520, 2838, 3338, -2996, -3148, 3134, 2983, -3273, 
-2839, 3396, 2688, -3507, -2574, 3609, 2464, -3695, -2375, 
3760, 2296, -3804, -2227, 3839, 2183, -3851, -2150, 3844, 
2130, -3822, -2128, 3795, 2137, -3744, -2155, 3661, 2194, 
-3572, -2232, 3472, 2286, -3352, -2342, 3222, 2413, -3077, 
-2491, 2919, 2564, -2733, -2643, 2561, 2735, -2366, -2814, 
2160, 2902, -1940, -2972, 1719, 3052, -1489, -3131, 1264, 
3204, -1015, -3255, 779, 3311, -538, -3360, 304, 3388, 
-66, -3411, -159, 3425, 394, -3437, -613, 3424, 836, 
-3404, -1057, 3362, 1260, -3312, -1451, 3261, 1629, -3179, 
-1792, 3100, 1958, -3001, -2092, 2898, 2217, -2776, -2342, 
2663, 2436, -2531, -2523, 2384, 2595, -2237, -2648, 2095, 
2684, -1929, -2703, 1768, 2704, -1611, -2685, 1452, 2655, 
-1298, -2608, 1128, 2555, -983, -2481, 823, 2391, -688, 
-2277, 550, 2157, -422, -2024, 294, 1874, -184, -1730, 
83, 1560, 2, -1373, -92, 1187, 154, -997, -205, 
781, 254, -573, -278, 356, 293, -140, -292, -89, 
276, 316, -249, -548, 206, 794, -158, -1015, 101, 
1255, -23, -1499, -65, 1728, 142, -1962, -257, 2177, 
354, -2413, -481, 2626, 585, -2852, -719, 3064, 847, 
-3259, -968, 3457, 1088, -3660, -1220, 3838, 1339, -4014, 
-1467, 4189, 1586, -4357, -1689, 4508, 1806, -4644, -1896, 
4784, 1980, -4925, -2067, 5038, 2123, -5154, -2183, 5245, 
2224, -5343, -2259, 5430, 2286, -5496, -2297, 5566, 2283, 
-5614, -2261, 5658, 2238, -5693, -2199, 5720, 2131, -5736, 
-2072, 5747, 1998, -5739, -1896, 5735, 1805, -5716, -1690, 
5685, 1585, -5646, -1459, 5596, 1323, -5539, -1186, 5467, 
1039, -5394, -899, 5319, 742, -5218, -596, 5129, 450, 
-5019, -301, 4905, 143, -4795, -8, 4663, -132, -4528, 
258, 4384, -394, -4242, 514, 4086, -634, -3938, 728, 
3776, -831, -3615, 915, 3435, -995, -3265, 1055, 3083, 
-1110, -2912, 1144, 2728, -1181, -2554, 1202, 2364, -1216, 
-2186, 1213, 2009, -1197, -1830, 1185, 1648, -1153, -1477, 
1109, 1289, -1053, -1130, 998, 964, -931, -809, 861, 
645, -802, -500, 716, 367, -644, -234, 554, 114, 
-465, 10, 387, -123, -309, 215, 222, -303, -147, 
377, 78, -455, -1, 503, -54, -547, 112, 589, 
-165, -624, 206, 638, -228, -630, 248, 627, -264, 
-614, 272, 586, -249, -556, 230, 507, -207, -440, 
165, 391, -116, -310, 42, 237, 17, -158, -103, 
69, 194, 39, -299, -134, 410, 228, -525, -338, 
659, 456, -779, -559, 927, 667, -1063, -775, 1206, 
879, -1350, -974, 1508, 1084, -1651, -1164, 1805, 1265, 
-1948, -1348, 2086, 1424, -2238, -1483, 2361, 1537, -2501, 
-1590, 2631, 1624, -2743, -1660, 2855, 1681, -2951, -1679, 
3056, 1689, -3126, -1670, 3196, 1640, -3268, -1596, 3325, 
1539, -3358, -1482, 3379, 1412, -3394, -1319, 3404, 1226, 
-3388, -1109, 3373, 988, -3343, -865, 3302, 729, -3250, 
-571, 3180, 418, -3113, -258, 3023, 93, -2928, 81, 
2817, -268, -2716, 447, 2593, -630, -2465, 825, 2340, 
-1014, -2200, 1198, 2057, -1378, -1907, 1569, 1768, -1755, 
-1620, 1935, 1461, -2094, -1313, 2275, 1154, -2424, -1009, 
2583, 850, -2727, -695, 2866, 556, -2992, -409, 3110, 
266, -3207, -141, 3298, -2, -3378, 124, 3460, -247, 
-3510, 352, 3561, -461, -3583, 563, 3607, -665, -3623, 
755, 3606, -836, -3597, 921, 3563, -996, -3528, 1047, 
3484, -1112, -3407, 1165, 3341, -1200, -3254, 1249, 3166, 
-1280, -3078, 1311, 2972, -1322, -2852, 1333, 2726, -1350, 
-2598, 1350, 2479, -1348, -2345, 1335, 2210, -1333, -2064, 
1316, 1927, -1295, -1786, 1256, 1636, -1239, -1500, 1201, 
1360, -1157, -1223, 1116, 1083, -1072, -944, 1020, 821, 
-964, -694, 900, 587, -826, -467, 760, 371, -694, 
-268, 611, 180, -534, -92, 446, 5, -362, 53, 
278, -129, -183, 178, 92, -230, 15, 278, -127, 
-301, 224, 336, -338, -349, 453, 364, -575, -361, 
693, 357, -812, -354, 937, 331, -1059, -307, 1180, 
290, -1316, -257, 1431, 204, -1571, -168, 1688, 118, 
-1824, -74, 1947, 12, -2075, 50, 2207, -108, -2325, 
163, 2438, -235, -2552, 306, 2658, -374, -2776, 454, 
2879, -524, -2981, 594, 3058, -670, -3155, 757, 3234, 
-832, -3303, 905, 3367, -982, -3433, 1052, 3471, -1126, 
-3517, 1206, 3564, -1271, -3588, 1343, 3608, -1421, -3618, 
1484, 3621, -1563, -3621, 1628, 3619, -1694, -3600, 1751, 
3578, -1815, -3542, 1868, 3504, -1929, -3463, 1986, 3402, 
-2037, -3352, 2074, 3303, -2123, -3239, 2162, 3169, -2214, 
-3112, 2245, 3031, -2268, -2967, 2291, 2901, -2317, -2819, 
2338, 2755, -2346, -2686, 2364, 2627, -2352, -2561, 2348, 
2495, -2348, -2440, 2335, 2379, -2307, -2334, 2283, 2297, 
-2245, -2255, 2191, 2217, -2155, -2189, 2088, 2168, -2035, 
-2147, 1952, 2134, -1873, -2136, 1790, 2134, -1699, -2125, 
1595, 2142, -1479, -2151, 1364, 2162, -1226, -2190, 1096, 
2212, -967, -2231, 809, 2261, -662, -2290, 493, 2311, 
-325, -2343, 155, 2372, 10, -2388, -200, 2407, 383, 
-2415, -563, 2420, 758, -2421, -957, 2419, 1154, -2411, 
-1342, 2379, 1549, -2353, -1742, 2306, 1932, -2252, -2128, 
2194, 2318, -2128, -2516, 2029, 2703, -1933, -2877, 1831, 
3059, -1707, -3227, 1572, 3393, -1412, -3539, 1261, 3692, 
-1082, -3827, 901, 3967, -710, -4083, 513, 4196, -294, 
-4300, 67, 4378, 154, -4464, -397, 4533, 634, -4583, 
-870, 4623, 1127, -4667, -1379, 4680, 1628, -4682, -1861, 
4690, 2113, -4672, -2343, 4644, 2582, -4600, -2809, 4553, 
3018, -4482, -3232, 4424, 3415, -4336, -3593, 4244, 3769, 
-4143, -3916, 4030, 4043, -3908, -4159, 3786, 4252, -3637, 
-4324, 3493, 4379, -3351, -4406, 3204, 4402, -3044, -4388, 
2868, 4347, -2705, -4292, 2530, 4195, -2364, -4097, 2183, 
3958, -2011, -3807, 1823, 3632, -1652, -3428, 1472, 3208, 
-1296, -2974, 1115, 2706, -935, -2440, 757, 2148, -586, 
-1843, 426, 1528, -262, -1200, 99, 860, 67, -530, 
-222, 177, 367, 178, -518, -523, 659, 888, -809, 
-1221, 933, 1580, -1076, -1916, 1192, 2249, -1319, -2565, 
1432, 2873, -1555, -3169, 1668, 3435, -1775, -3707, 1876, 
3954, -1973, -4177, 2066, 4378, -2156, -4554, 2245, 4714, 
-2329, -4853, 2421, 4961, -2496, -5038, 2574, 5114, -2645, 
-5141, 2718, 5152, -2780, -5131, 2847, 5107, -2908, -5031, 
2971, 4957, -3041, -4841, 3092, 4718, -3154, -4566, 3197, 
4391, -3250, -4193, 3296, 3992, -3336, -3767, 3387, 3541, 
-3432, -3291, 3475, 3022, -3510, -2751, 3539, 2493, -3561, 
-2209, 3588, 1915, -3623, -1635, 3644, 1354, -3654, -1074, 
3678, 795, -3682, -510, 3698, 248, -3702, 23, 3700, 
-273, -3698, 501, 3690, -737, -3682, 943, 3667, -1143, 
-3648, 1342, 3626, -1510, -3600, 1654, 3587, -1794, -3556, 
1915, 3518, -2012, -3482, 2093, 3435, -2162, -3388, 2211, 
3342, -2254, -3289, 2268, 3229, -2265, -3178, 2240, 3119, 
-2222, -3045, 2176, 2986, -2108, -2920, 2039, 2853, -1968, 
-2767, 1876, 2701, -1771, -2630, 1676, 2553, -1570, -2470, 
1453, 2402, -1329, -2317, 1211, 2237, -1079, -2166, 967, 
2079, -840, -2007, 728, 1922, -620, -1844, 510, 1760, 
-406, -1695, 305, 1614, -225, -1529, 152, 1461, -79, 
-1387, 14, 1317, 31, -1237, -73, 1173, 96, -1100, 
-106, 1030, 114, -972, -119, 908, 91, -837, -73, 
784, 30, -715, 23, 675, -73, -606, 147, 557, 
-218, -522, 298, 465, -387, -421, 478, 397, -584, 
-359, 699, 326, -803, -301, 919, 277, -1036, -255, 
1142, 239, -1254, -219, 1380, 213, -1488, -207, 1598, 
221, -1704, -226, 1810, 238, -1892, -260, 1984, 285, 
-2071, -324, 2157, 364, -2215, -411, 2273, 455, -2334, 
-511, 2383, 574, -2411, -654, 2448, 730, -2468, -806, 
2471, 902, -2475, -1008, 2474, 1110, -2445, -1216, 2425, 
1326, -2393, -1453, 2351, 1580, -2316, -1708, 2255, 1831, 
-2214, -1972, 2150, 2115, -2088, -2249, 2019, 2399, -1941, 
-2548, 1868, 2685, -1797, -2825, 1727, 2961, -1647, -3116, 
1588, 3247, -1518, -3382, 1438, 3509, -1383, -3629, 1316, 
3741, -1275, -3839, 1213, 3945, -1185, -4034, 1151, 4113, 
-1115, -4178, 1096, 4235, -1075, -4286, 1071, 4313, -1077, 
-4318, 1097, 4330, -1111, -4317, 1145, 4287, -1179, -4237, 
1230, 4187, -1283, -4105, 1341, 4008, -1414, -3904, 1502, 
3783, -1593, -3650, 1683, 3497, -1788, -3314, 1891, 3141, 
-2003, -2949, 2125, 2744, -2237, -2516, 2375, 2290, -2491, 
-2046, 2627, 1801, -2755, -1542, 2900, 1290, -3036, -1023, 
3171, 755, -3302, -480, 3432, 202, -3575, 51, 3698, 
-315, -3831, 575, 3940, -842, -4066, 1073, 4184, -1312, 
-4281, 1543, 4394, -1744, -4479, 1951, 4581, -2125, -4661, 
2284, 4735, -2430, -4815, 2562, 4870, -2667, -4932, 2752, 
4980, -2813, -5028, 2836, 5062, -2862, -5087, 2848, 5108, 
-2819, -5115, 2756, 5121, -2666, -5120, 2569, 5117, -2429, 
-5098, 2276, 5069, -2108, -5055, 1914, 5026, -1692, -4983, 
1449, 4950, -1199, -4902, 915, 4859, -620, -4810, 320, 
4763, -7, -4707, -319, 4645, 644, -4595, -997, 4542, 
1338, -4476, -1695, 4426, 2039, -4363, -2376, 4307, 2731, 
-4254, -3070, 4215, 3395, -4165, -3720, 4114, 4024, -4080, 
-4312, 4030, 4591, -4010, -4848, 3974, 5090, -3955, -5303, 
3926, 5511, -3917, -5680, 3910, 5823, -3901, -5949, 3896, 
6054, -3898, -6118, 3920, 6152, -3934, -6169, 3947, 6167, 
-3977, -6127, 4016, 6054, -4049, -5950, 4100, 5828, -4145, 
-5691, 4196, 5522, -4242, -5324, 4299, 5099, -4374, -4864, 
4437, 4607, -4502, -4331, 4570, 4040, -4638, -3723, 4714, 
3407, -4787, -3090, 4857, 2739, -4928, -2407, 4991, 2063, 
-5054, -1705, 5133, 1358, -5191, -1022, 5254, 673, -5305, 
-349, 5348, 30, -5397, 289, 5429, -590, -5471, 866, 
5496, -1142, -5513, 1403, 5511, -1637, -5519, 1837, 5521, 
-2035, -5500, 2214, 5462, -2359, -5439, 2478, 5389, -2581, 
-5326, 2653, 5259, -2708, -5181, 2744, 5100, -2750, -5008, 
2724, 4896, -2679, -4779, 2628, 4646, -2549, -4498, 2444, 
4358, -2313, -4198, 2168, 4037, -2023, -3848, 1858, 3673, 
-1661, -3482, 1470, 3281, -1265, -3079, 1069, 2869, -837, 
-2654, 630, 2443, -394, -2220, 184, 1989, 40, -1760, 
-260, 1548, 479, -1320, -685, 1101, 886, -871, -1077, 
654, 1246, -436, -1413, 223, 1563, -31, -1711, -173, 
1822, 371, -1923, -543, 2022, 716, -2083, -897, 2146, 
1046, -2180, -1191, 2185, 1334, -2179, -1447, 2157, 1563, 
-2112, -1673, 2055, 1749, -1992, -1825, 1889, 1894, -1794, 
-1956, 1670, 2000, -1530, -2019, 1388, 2052, -1229, -2056, 
1046, 2055, -876, -2038, 688, 2023, -499, -1977, 294, 
1948, -97, -1902, -98, 1844, 306, -1794, -498, 1721, 
707, -1650, -899, 1588, 1090, -1515, -1266, 1429, 1454, 
-1355, -1611, 1277, 1768, -1207, -1920, 1138, 2050, -1058, 
-2179, 994, 2291, -939, -2396, 894, 2478, -835, -2555, 
797, 2614, -772, -2653, 741, 2681, -725, -2702, 708, 
2714, -719, -2700, 730, 2673, -744, -2653, 771, 2606, 
-805, -2541, 855, 2480, -924, -2407, 982, 2326, -1057, 
-2236, 1134, 2140, -1234, -2040, 1318, 1931, -1432, -1816, 
1542, 1700, -1648, -1583, 1763, 1476, -1879, -1362, 2009, 
1246, -2133, -1129, 2252, 1023, -2364, -918, 2487, 826, 
-2603, -728, 2724, 641, -2824, -546, 2937, 474, -3024, 
-413, 3112, 351, -3197, -287, 3255, 239, -3326, -207, 
3371, 188, -3421, -166, 3440, 144, -3464, -137, 3456, 
146, -3458, -156, 3437, 171, -3399, -206, 3359, 242, 
-3308, -280, 3233, 315, -3148, -362, 3064, 426, -2966, 
-486, 2849, 536, -2737, -603, 2602, 670, -2468, -746, 
2322, 822, -2174, -889, 2028, 951, -1871, -1035, 1703, 
1103, -1557, -1170, 1395, 1249, -1225, -1314, 1077, 1381, 
-919, -1437, 771, 1506, -636, -1564, 490, 1610, -376, 
-1669, 246, 1716, -140, -1755, 35, 1795, 42, -1844, 
-119, 1873, 190, -1907, -233, 1929, 276, -1951, -305, 
1958, 303, -1977, -312, 1991, 285, -1992, -250, 2005, 
205, -2008, -140, 1994, 68, -1991, 23, 1974, -118, 
-1967, 232, 1949, -353, -1934, 491, 1900, -637, -1884, 
788, 1854, -947, -1812, 1120, 1779, -1299, -1729, 1472, 
1680, -1663, -1632, 1853, 1589, -2046, -1525, 2232, 1470, 
-2413, -1397, 2607, 1341, -2793, -1271, 2972, 1181, -3151, 
-1104, 3327, 1027, -3503, -936, 3654, 838, -3807, -736, 
3968, 637, -4107, -524, 4222, 422, -4348, -305, 4461, 
192, -4559, -71, 4645, -52, -4713, 175, 4787, -310, 
-4839, 435, 4879, -554, -4913, 681, 4948, -808, -4952, 
947, 4962, -1068, -4956, 1194, 4949, -1319, -4925, 1431, 
4898, -1547, -4860, 1655, 4809, -1745, -4768, 1849, 4707, 
-1931, -4650, 2005, 4590, -2071, -4509, 2126, 4449, -2181, 
-4371, 2219, 4301, -2247, -4226, 2256, 4142, -2257, -4077, 
2243, 3989, -2220, -3914, 2176, 3834, -2120, -3767, 2061, 
3687, -1970, -3612, 1877, 3535, -1770, -3469, 1634, 3398, 
-1502, -3328, 1357, 3260, -1188, -3183, 1029, 3126, -836, 
-3050, 638, 2992, -445, -2918, 228, 2853, -22, -2775, 
-204, 2714, 429, -2635, -658, 2576, 898, -2487, -1117, 
2410, 1355, -2335, -1583, 2240, 1814, -2148, -2021, 2058, 
2244, -1962, -2446, 1862, 2641, -1744, -2816, 1643, 2992, 
-1527, -3153, 1398, 3301, -1277, -3420, 1141, 3540, -1013, 
-3620, 865, 3704, -717, -3761, 576, 3801, -421, -3809, 
270, 3806, -113, -3800, -57, 3757, 209, -3686, -363, 
3607, 529, -3504, -697, 3378, 846, -3252, -1001, 3090, 
1168, -2915, -1306, 2731, 1462, -2518, -1597, 2307, 1741, 
-2086, -1868, 1848, 1980, -1600, -2092, 1333, 2208, -1078, 
-2303, 810, 2390, -546, -2471, 275, 2529, 1, -2597, 
-255, 2638, 526, -2676, -775, 2694, 1026, -2719, -1264, 
2711, 1499, -2713, -1726, 2703, 1936, -2675, -2132, 2629, 
2311, -2590, -2467, 2534, 2608, -2483, -2747, 2419, 2860, 
-2350, -2960, 2262, 3034, -2188, -3087, 2103, 3123, -2011, 
-3157, 1921, 3149, -1837, -3136, 1739, 3119, -1657, -3074, 
1562, 3002, -1487, -2929, 1407, 2843, -1341, -2750, 1268, 
2625, -1216, -2516, 1158, 2380, -1129, -2253, 1095, 2107, 
-1066, -1960, 1048, 1823, -1062, -1665, 1063, 1521, -1085, 
-1376, 1125, 1233, -1168, -1097, 1226, 962, -1298, -833, 
1389, 721, -1475, -626, 1583, 525, -1703, -444, 1831, 
369, -1967, -295, 2108, 250, -2263, -209, 2414, 185, 
-2575, -187, 2758, 185, -2931, -200, 3108, 233, -3283, 
-275, 3454, 328, -3639, -383, 3805, 457, -3988, -536, 
4161, 616, -4320, -715, 4471, 816, -4633, -910, 4780, 
1017, -4911, -1120, 5035, 1230, -5137, -1337, 5244, 1443, 
-5340, -1529, 5404, 1630, -5474, -1716, 5520, 1793, -5559, 
-1850, 5572, 1901, -5581, -1946, 5565, 1978, -5541, -2001, 
5513, 2012, -5457, -2000, 5393, 1971, -5313, -1933, 5207, 
1873, -5110, -1803, 4982, 1724, -4854, -1616, 4727, 1490, 
-4576, -1359, 4420, 1227, -4255, -1071, 4085, 902, -3906, 
-717, 3720, 519, -3528, -333, 3348, 120, -3151, 77, 
2965, -295, -2769, 512, 2590, -720, -2403, 936, 2212, 
-1145, -2029, 1350, 1855, -1550, -1690, 1754, 1527, -1925, 
-1360, 2101, 1214, -2261, -1068, 2405, 947, -2538, -811, 
2652, 701, -2754, -603, 2818, 496, -2885, -413, 2925, 
333, -2947, -273, 2945, 218, -2914, -163, 2880, 123, 
-2814, -96, 2721, 73, -2614, -63, 2488, 50, -2353, 
-49, 2193, 72, -2015, -72, 1813, 109, -1605, -128, 
1395, 165, -1160, -202, 919, 250, -674, -286, 413, 
347, -149, -390, -98, 442, 368, -499, -628, 553, 
878, -622, -1128, 678, 1377, -745, -1605, 802, 1822, 
-870, -2038, 920, 2224, -977, -2412, 1041, 2567, -1108, 
-2700, 1164, 2835, -1220, -2929, 1267, 3010, -1333, -3065, 
1383, 3103, -1437, -3121, 1483, 3112, -1520, -3075, 1573, 
3015, -1624, -2925, 1667, 2823, -1702, -2696, 1751, 2552, 
-1774, -2384, 1816, 2193, -1847, -1987, 1888, 1765, -1903, 
-1524, 1936, 1277, -1968, -1007, 1988, 744, -2003, -450, 
2011, 168, -2026, 126, 2034, -419, -2037, 721, 2028, 
-1026, -2026, 1333, 2026, -1618, -2008, 1918, 1978, -2202, 
-1957, 2467, 1913, -2725, -1872, 2980, 1836, -3229, -1775, 
3449, 1714, -3660, -1650, 3864, 1567, -4046, -1490, 4194, 
1404, -4343, -1297, 4471, 1199, -4570, -1086, 4671, 967, 
-4742, -826, 4793, 699, -4817, -568, 4838, 420, -4842, 
-265, 4823, 107, -4790, 43, 4728, -216, -4679, 371, 
4604, -540, -4506, 705, 4403, -862, -4297, 1039, 4188, 
-1204, -4060, 1357, 3917, -1503, -3794, 1666, 3646, -1803, 
-3501, 1943, 3360, -2060, -3210, 2187, 3051, -2289, -2918, 
2374, 2764, -2456, -2613, 2522, 2480, -2585, -2345, 2627, 
2205, -2645, -2082, 2646, 1960, -2631, -1838, 2601, 1724, 
-2568, -1621, 2491, 1507, -2421, -1419, 2317, 1317, -2207, 
-1227, 2057, 1148, -1909, -1053, 1744, 973, -1570, -901, 
1363, 824, -1153, -741, 938, 671, -694, -586, 446, 
506, -203, -423, -70, 337, 327, -251, -603, 166, 
887, -60, -1160, -38, 1429, 148, -1707, -253, 1972, 
383, -2237, -512, 2495, 647, -2723, -792, 2958, 942, 
-3184, -1099, 3390, 1266, -3572, -1433, 3743, 1618, -3883, 
-1801, 4016, 1981, -4136, -2173, 4213, 2371, -4269, -2586, 
4323, 2785, -4336, -3001, 4324, 3200, -4274, -3406, 4221, 
3618, -4133, -3817, 4031, 4032, -3890, -4220, 3728, 4417, 
-3550, -4598, 3347, 4784, -3125, -4948, 2875, 5113, -2609, 
-5259, 2344, 5401, -2041, -5523, 1741, 5624, -1419, -5727, 
1100, 5810, -759, -5887, 434, 5927, -83, -5976, -258, 
5996, 589, -5997, -935, 5981, 1266, -5951, -1579, 5913, 
1891, -5838, -2207, 5772, 2493, -5677, -2762, 5575, 3020, 
-5446, -3264, 5324, 3471, -5171, -3679, 5024, 3849, -4851, 
-4007, 4680, 4126, -4487, -4228, 4298, 4322, -4105, -4375, 
3910, 4408, -3700, -4414, 3484, 4381, -3282, -4354, 3072, 
4278, -2866, -4200, 2649, 4088, -2452, -3961, 2255, 3810, 
-2056, -3655, 1866, 3476, -1684, -3278, 1514, 3068, -1343, 
-2868, 1180, 2641, -1030, -2411, 889, 2170, -742, -1946, 
626, 1706, -513, -1468, 407, 1238, -309, -1014, 229, 
793, -137, -590, 65, 396, 0, -210, -43, 26, 
99, 126, -147, -263, 185, 400, -212, -501, 246, 
593, -258, -669, 280, 726, -308, -750, 321, 776, 
-346, -769, 364, 746, -384, -716, 393, 665, -414, 
-592, 443, 517, -467, -412, 490, 305, -533, -188, 
555, 63, -595, 70, 626, -199, -673, 336, 714, 
-490, -769, 625, 803, -761, -866, 899, 916, -1014, 
-952, 1138, 1009, -1258, -1053, 1347, 1102, -1436, -1146, 
1507, 1196, -1560, -1224, 1603, 1263, -1615, -1289, 1622, 
1311, -1599, -1312, 1561, 1316, -1498, -1305, 1424, 1303, 
-1330, -1273, 1211, 1243, -1064, -1191, 902, 1134, -728, 
-1064, 541, 980, -326, -885, 93, 782, 151, -667, 
-392, 529, 656, -401, -940, 245, 1222, -82, -1505, 
-73, 1778, 253, -2074, -442, 2347, 633, -2635, -821, 
2908, 1021, -3162, -1223, 3429, 1429, -3670, -1627, 3892, 
1828, -4103, -2024, 4295, 2216, -4465, -2397, 4610, 2574, 
-4730, -2729, 4838, 2885, -4918, -3023, 4964, 3142, -4989, 
-3240, 4968, 3342, -4937, -3405, 4880, 3464, -4789, -3485, 
4670, 3494, -4538, -3479, 4359, 3442, -4175, -3377, 3952, 
3300, -3713, -3202, 3454, 3059, -3167, -2917, 2882, 2741, 
-2560, -2541, 2250, 2313, -1909, -2079, 1580, 1818, -1227, 
-1541, 883, 1258, -544, -962, 188, 643, 151, -310, 
-470, -15, 788, 364, -1101, -702, 1381, 1048, -1664, 
-1394, 1920, 1748, -2139, -2076, 2351, 2407, -2521, -2736, 
2682, 3046, -2807, -3337, 2895, 3613, -2954, -3857, 2988, 
4091, -2986, -4309, 2947, 4494, -2876, -4659, 2769, 4790, 
-2651, -4879, 2472, 4957, -2288, -5008, 2061, 5010, -1809, 
-4994, 1541, 4939, -1230, -4845, 906, 4740, -557, -4584, 
192, 4416, 185, -4199, -570, 3971, 983, -3703, -1389, 
3417, 1803, -3109, -2233, 2772, 2658, -2419, -3066, 2052, 
3474, -1672, -3884, 1273, 4268, -864, -4655, 461, 5018, 
-47, -5357, -381, 5678, 788, -5968, -1203, 6251, 1601, 
-6491, -1994, 6715, 2372, -6897, -2728, 7052, 3079, -7177, 
-3395, 7275, 3704, -7337, -3977, 7357, 4221, -7356, -4438, 
7306, 4631, -7237, -4795, 7135, 4908, -6994, -5001, 6835, 
5066, -6633, -5088, 6403, 5079, -6152, -5027, 5879, 4950, 
-5592, -4834, 5274, 4680, -4944, -4503, 4595, 4289, -4227, 
-4057, 3843, 3777, -3471, -3487, 3067, 3182, -2676, -2841, 
2284, 2479, -1890, -2122, 1500, 1731, -1108, -1339, 735, 
928, -372, -524, 18, 107, 330, 295, -654, -700, 
971, 1092, -1258, -1485, 1529, 1872, -1784, -2235, 2006, 
2585, -2225, -2912, 2402, 3221, -2569, -3500, 2706, 3765, 
-2819, -3996, 2903, 4193, -2969, -4368, 3024, 4506, -3051, 
-4629, 3057, 4698, -3040, -4751, 2993, 4765, -2952, -4748, 
2887, 4713, -2804, -4631, 2701, 4526, -2600, -4394, 2491, 
4226, -2365, -4042, 2229, 3830, -2097, -3583, 1957, 3333, 
-1820, -3049, 1670, 2765, -1547, -2459, 1405, 2148, -1279, 
-1810, 1157, 1484, -1040, -1147, 934, 811, -835, -471, 
751, 142, -668, 193, 600, -506, -550, 819, 506, 
-1107, -476, 1394, 474, -1664, -462, 1913, 477, -2139, 
-487, 2339, 536, -2523, -573, 2689, 628, -2814, -698, 
2929, 762, -3008, -845, 3074, 930, -3114, -1031, 3108, 
1122, -3102, -1218, 3065, 1332, -2994, -1430, 2907, 1527, 
-2795, -1630, 2660, 1733, -2512, -1816, 2344, 1916, -2166, 
-1996, 1964, 2073, -1765, -2139, 1538, 2191, -1302, -2235, 
1078, 2280, -832, -2313, 587, 2322, -355, -2332, 111, 
2308, 136, -2295, -367, 2264, 592, -2226, -797, 2168, 
1013, -2099, -1203, 2023, 1377, -1943, -1553, 1835, 1695, 
-1740, -1838, 1628, 1956, -1517, -2039, 1392, 2131, -1260, 
-2181, 1138, 2229, -1001, -2239, 873, 2253, -736, -2231, 
613, 2203, -483, -2145, 361, 2083, -237, -1992, 121, 
1892, -19, -1775, -65, 1654, 161, -1516, -221, 1364, 
293, -1216, -339, 1047, 385, -883, -413, 715, 427, 
-545, -413, 383, 406, -201, -370, 45, 340, 115, 
-282, -269, 210, 413, -130, -552, 45, 678, 73, 
-809, -181, 900, 298, -1003, -444, 1075, 583, -1134, 
-727, 1182, 880, -1202, -1027, 1221, 1185, -1211, -1357, 
1190, 1507, -1157, -1671, 1108, 1820, -1027, -1985, 943, 
2127, -847, -2265, 724, 2400, -594, -2519, 462, 2640, 
-310, -2745, 143, 2834, 34, -2913, -216, 2978, 405, 
-3021, -588, 3063, 789, -3081, -992, 3084, 1189, -3074, 
-1400, 3055, 1602, -3004, -1808, 2946, 2005, -2881, -2196, 
2798, 2381, -2699, -2548, 2583, 2718, -2467, -2890, 2324, 
3027, -2174, -3176, 2028, 3300, -1871, -3414, 1697, 3517, 
-1530, -3614, 1358, 3680, -1168, -3743, 991, 3801, -823, 
-3823, 645, 3853, -469, -3861, 297, 3861, -149, -3838, 
-14, 3804, 153, -3767, -284, 3713, 388, -3641, -491, 
3568, 582, -3500, -652, 3408, 713, -3311, -761, 3207, 
776, -3095, -779, 2990, 770, -2883, -725, 2763, 678, 
-2651, -601, 2532, 493, -2423, -389, 2311, 247, -2205, 
-107, 2088, -72, -1993, 250, 1903, -468, -1810, 681, 
1729, -920, -1657, 1161, 1586, -1414, -1521, 1697, 1476, 
-1969, -1433, 2257, 1404, -2551, -1395, 2847, 1386, -3146, 
-1377, 3446, 1392, -3753, -1401, 4060, 1428, -4355, -1471, 
4652, 1511, -4926, -1574, 5220, 1639, -5480, -1715, 5749, 
1790, -5990, -1877, 6217, 1965, -6445, -2056, 6651, 2163, 
-6840, -2278, 7004, 2376, -7159, -2505, 7295, 2621, -7414, 
-2743, 7505, 2851, -7575, -2980, 7630, 3092, -7657, -3226, 
7676, 3340, -7679, -3455, 7652, 3568, -7601, -3687, 7539, 
3783, -7440, -3895, 7342, 4001, -7223, -4095, 7079, 4180, 
-6937, -4264, 6760, 4346, -6583, -4413, 6379, 4477, -6178, 
-4537, 5961, 4575, -5732, -4622, 5482, 4652, -5245, -4670, 
4987, 4699, -4738, -4707, 4467, 4707, -4200, -4685, 3929, 
4672, -3676, -4648, 3398, 4608, -3136, -4577, 2873, 4518, 
-2617, -4452, 2351, 4386, -2105, -4306, 1851, 4212, -1615, 
-4113, 1367, 4018, -1141, -3903, 925, 3784, -720, -3651, 
506, 3507, -314, -3368, 133, 3220, 46, -3054, -211, 
2882, 369, -2706, -525, 2533, 658, -2351, -796, 2155, 
912, -1961, -1030, 1749, 1129, -1551, -1217, 1344, 1296, 
-1127, -1371, 903, 1452, -688, -1503, 461, 1561, -242, 
-1603, 16, 1633, 204, -1654, -419, 1676, 649, -1702, 
-871, 1712, 1082, -1713, -1301, 1706, 1516, -1697, -1733, 
1669, 1927, -1647, -2129, 1616, 2327, -1579, -2513, 1546, 
2685, -1490, -2850, 1437, 3027, -1379, -3168, 1315, 3326, 
-1253, -3458, 1167, 3588, -1093, -3703, 998, 3803, -898, 
-3894, 804, 3978, -693, -4046, 585, 4113, -470, -4169, 
342, 4201, -225, -4235, 90, 4251, 59, -4251, -200, 
4257, 343, -4233, -512, 4207, 663, -4184, -822, 4136, 
988, -4080, -1162, 4032, 1339, -3969, -1522, 3898, 1696, 
-3822, -1874, 3739, 2046, -3649, -2236, 3556, 2423, -3454, 
-2593, 3364, 2775, -3273, -2946, 3172, 3130, -3070, -3293, 
2975, 3455, -2880, -3621, 2795, 3769, -2698, -3905, 2625, 
4048, -2534, -4184, 2461, 4303, -2383, -4414, 2318, 4514, 
-2265, -4597, 2206, 4686, -2158, -4739, 2113, 4799, -2069, 
-4838, 2036, 4874, -2000, -4879, 1985, 4879, -1969, -4866, 
1955, 4850, -1956, -4809, 1948, 4761, -1940, -4694, 1948, 
4606, -1949, -4517, 1963, 4420, -1965, -4290, 1962, 4172, 
-1971, -4028, 1971, 3883, -1979, -3738, 1976, 3579, -1970, 
-3408, 1948, 3231, -1936, -3055, 1908, 2870, -1874, -2680, 
1834, 2485, -1780, -2299, 1715, 2108, -1635, -1925, 1552, 
1751, -1447, -1569, 1345, 1399, -1214, -1236, 1080, 1072, 
-938, -921, 775, 791, -600, -648, 416, 538, -219, 
-433, 21, 332, 203, -269, -442, 194, 682, -141, 
-934, 111, 1201, -96, -1460, 91, 1734, -103, -2014, 
118, 2308, -159, -2601, 214, 2880, -284, -3181, 382, 
3462, -467, -3756, 580, 4041, -709, -4320, 830, 4606, 
-978, -4874, 1125, 5129, -1286, -5379, 1449, 5619, -1619, 
-5836, 1792, 6052, -1968, -6240, 2134, 6425, -2317, -6582, 
2498, 6734, -2660, -6856, 2825, 6961, -2987, -7042, 3132, 
7115, -3280, -7148, 3422, 7171, -3527, -7169, 3644, 7152, 
-3744, -7123, 3824, 7065, -3887, -6981, 3931, 6875, -3956, 
-6756, 3966, 6621, -3963, -6465, 3939, 6294, -3879, -6108, 
3814, 5898, -3734, -5693, 3637, 5459, -3514, -5228, 3366, 
4974, -3204, -4725, 3016, 4462, -2815, -4202, 2609, 3924, 
-2377, -3662, 2133, 3386, -1881, -3124, 1612, 2850, -1334, 
-2592, 1038, 2333, -739, -2090, 434, 1864, -116, -1629, 
-184, 1413, 499, -1215, -820, 1017, 1138, -844, -1438, 
682, 1747, -525, -2043, 402, 2341, -284, -2624, 194, 
2892, -114, -3141, 53, 3381, 0, -3620, -21, 3824, 
33, -4020, -29, 4202, 18, -4357, 15, 4494, -61, 
-4598, 138, 4698, -198, -4765, 294, 4827, -385, -4855, 
489, 4868, -606, -4854, 739, 4822, -868, -4762, 994, 
4676, -1128, -4590, 1275, 4469, -1406, -4350, 1552, 4200, 
-1689, -4030, 1815, 3854, -1936, -3656, 2070, 3464, -2174, 
-3249, 2276, 3030, -2378, -2794, 2464, 2551, -2535, -2313, 
2610, 2071, -2654, -1823, 2697, 1575, -2720, -1330, 2724, 
1093, -2730, -867, 2707, 625, -2675, -412, 2612, 186, 
-2558, 4, 2479, -197, -2380, 382, 2269, -549, -2156, 
712, 2008, -850, -1863, 965, 1709, -1074, -1540, 1165, 
1351, -1248, -1171, 1310, 976, -1355, -760, 1368, 557, 
-1379, -331, 1369, 116, -1350, 111, 1321, -323, -1268, 
552, 1201, -776, -1115, 1001, 1025, -1212, -925, 1430, 
807, -1649, -692, 1854, 559, -2050, -408, 2242, 262, 
-2416, -109, 2582, -45, -2751, 199, 2900, -369, -3030, 
520, 3147, -681, -3266, 844, 3358, -1009, -3450, 1157, 
3513, -1321, -3565, 1464, 3600, -1611, -3632, 1732, 3645, 
-1869, -3641, 1987, 3620, -2103, -3581, 2192, 3544, -2289, 
-3476, 2377, 3410, -2454, -3322, 2510, 3220, -2579, -3106, 
2620, 2997, -2652, -2853, 2688, 2719, -2694, -2565, 2707, 
2410, -2717, -2238, 2702, 2081, -2700, -1901, 2675, 1707, 
-2659, -1522, 2624, 1338, -2584, -1156, 2552, 949, -2503, 
-768
		)
		)
 port map ( 
			Clk_96 => Clk_96,
			Ce_F6 => Ce_F6,
			Sign_LCHM => Sign_LCHM,
			EN =>EN,
			Rom_cos_all => Rom_cos_L3_plus--out
			 );
----------------------------------


--------------------------------L40 ������ '-'
--LHM_PP1: entity work.LHM_ALL
--generic map(
--
--		rom_cos =>(8190, -302, -8161, 1102, 8052, -1892, -7868, 2663, 7605, -3410, -7272, 4121, 6867, -4795, -6399, 5421, 5866, -5997, -5280, 6513, 4642, -6968, -3961, 7355, 3240, -7673, -2490, 7915, 1715, -8084, 
---925, 8174, 125, -8187, 674, 8120, -1468, -7978, 2247, 7757, -3005, -7465, 3733, 7099, -4427, -6668, 5077, 6172, -5680, -5618, 6227, 5010, -6717, -4356, 7140, 3659, -7498, -2929, 7783, 2170, 
---7995, -1392, 8130, 599, -8189, 197, 8169, -993, -8073, 1778, 7899, -2547, -7652, 3291, 7331, -4005, -6943, 4679, 6487, -5310, -5972, 5890, 5399, -6415, -4777, 6878, 4108, -7278, -3402, 7607, 
--2663, -7867, -1900, 8050, 1118, -8159, -328, 8190, -467, -8146, 1256, 8023, -2035, -7827, 2792, 7555, -3525, -7215, 4223, 6805, -4883, -6333, 5495, 5801, -6057, -5216, 6561, 4580, -7005, -3903, 
--7381, 3189, -7691, -2446, 7926, 1679, -8089, -899, 8175, 108, -8186, 682, 8120, -1467, -7979, 2236, 7762, -2986, -7475, 3706, 7117, -4393, -6694, 5038, 6207, -5637, -5665, 6182, 5068, -6672, 
---4426, 7097, 3742, -7458, -3024, 7749, 2277, -7969, -1511, 8113, 730, -8185, 57, 8178, -844, -8098, 1622, 7941, -2386, -7713, 3126, 7411, -3839, -7043, 4515, 6609, -5151, -6115, 5737, 5563, 
---6272, -4963, 6747, 4314, -7162, -3628, 7509, 2907, -7789, -2161, 7995, 1394, -8129, -616, 8187, -169, -8172, 951, 8080, -1726, -7916, 2483, 7677, -3218, -7370, 3923, 6994, -4593, -6556, 5219, 
--6056, -5799, -5502, 6324, 4897, -6793, -4249, 7198, 3560, -7539, -2841, 7809, 2095, -8010, -1331, 8136, 554, -8190, 227, 8167, -1007, -8072, 1775, 7902, -2530, -7662, 3259, 7350, -3960, -6974, 
--4624, 6532, -5247, -6034, 5820, 5479, -6343, -4876, 6806, 4227, -7209, -3543, 7545, 2824, -7815, -2082, 8012, 1319, -8138, -547, 8189, -232, -8168, 1007, 8071, -1774, -7904, 2524, 7663, -3252, 
---7356, 3949, 6980, -4612, -6543, 5232, 6046, -5806, -5497, 6326, 4896, -6791, -4254, 7193, 3571, -7533, -2859, 7802, 2119, -8004, -1362, 8132, 592, -8189, 182, 8171, -956, -8081, 1719, 7918, 
---2469, -7685, 3194, 7382, -3893, -7016, 4554, 6584, -5177, -6097, 5752, 5553, -6277, -4961, 6744, 4324, -7153, -3650, 7497, 2942, -7775, -2210, 7982, 1456, -8121, -692, 8185, -80, -8178, 850, 
--8097, -1613, -7946, 2360, 7723, -3088, -7434, 3787, 7076, -4453, -6658, 5079, 6180, -5661, -5649, 6191, 5066, -6668, -4440, 7084, 3774, -7439, -3076, 7727, 2350, -7949, -1604, 8098, 843, -8179, 
---77, 8185, -692, -8121, 1452, 7984, -2202, -7778, 2930, 7503, -3634, -7163, 4304, 6759, -4938, -6298, 5526, 5780, -6068, -5213, 6555, 4598, -6986, -3946, 7354, 3257, -7660, -2542, 7897, 1803, 
---8066, -1050, 8163, 286, -8191, 478, 8145, -1239, -8031, 1988, 7844, -2721, -7591, 3428, 7270, -4108, -6888, 4749, 6444, -5351, -5947, 5904, 5395, -6408, -4799, 6854, 4160, -7242, -3486, 7566, 
--2781, -7826, -2054, 8016, 1307, -8139, -551, 8189, -212, -8170, 971, 8079, -1723, -7920, 2458, 7690, -3173, -7397, 3859, 7037, -4514, -6619, 5127, 6142, -5698, -5614, 6218, 5036, -6686, -4417, 
--7095, 3758, -7445, -3069, 7728, 2352, -7947, -1617, 8096, 866, -8177, -110, 8186, -649, -8127, 1401, 7996, -2142, -7799, 2862, 7533, -3560, -7205, 4225, 6814, -4856, -6366, 5443, 5862, -5986, 
---5310, 6475, 4711, -6911, -4074, 7286, 3400, -7601, -2700, 7849, 1975, -8032, -1235, 8145, 483, -8191, 271, 8165, -1025, -8071, 1768, 7907, -2497, -7679, 3203, 7383, -3884, -7026, 4530, 6608, 
---5139, -6136, 5702, 5611, -6219, -5040, 6682, 4425, -7089, -3774, 7435, 3090, -7720, -2382, 7938, 1652, -8091, -910, 8173, 159, -8189, 592, 8133, -1339, -8012, 2073, 7820, -2791, -7566, 3483, 
--7245, -4148, -6866, 4776, 6428, -5366, -5937, 5909, 5395, -6404, -4810, 6843, 4183, -7227, -3523, 7548, 2831, -7808, -2118, 8001, 1386, -8128, -644, 8186, -105, -8178, 851, 8099, -1592, -7954, 
--2317, 7742, -3024, -7467, 3705, 7128, -4356, -6732, 4969, 6277, -5542, -5773, 6068, 5219, -6544, -4624, 6964, 3988, -7329, -3322, 7630, 2626, -7870, -1911, 8043, 1178, -8151, -438, 8190, -308, 
---8163, 1050, 8067, -1784, -7906, 2501, 7677, -3200, -7388, 3870, 7035, -4510, -6627, 5110, 6162, -5671, -5648, 6182, 5087, -6644, -4485, 7050, 3845, -7400, -3175, 7686, 2477, -7912, -1761, 8071, 
--1029, -8165, -291, 8190, -451, -8150, 1188, 8042, -1917, -7869, 2627, 7631, -3319, -7332, 3980, 6971, -4611, -6555, 5203, 6084, -5753, -5565, 6255, 5000, -6707, -4395, 7103, 3753, -7443, -3083, 
--7720, 2385, -7936, -1670, 8086, 940, -8171, -205, 8189, -534, -8142, 1266, 8027, -1990, -7849, 2696, 7605, -3381, -7302, 4037, 6937, -4663, -6519, 5248, 6046, -5792, -5526, 6288, 4960, -6735, 
---4356, 7125, 3715, -7460, -3046, 7732, 2350, -7944, -1638, 8090, 911, -8173, -179, 8188, -556, -8139, 1285, 8023, -2005, -7845, 2707, 7601, -3389, -7298, 4042, 6935, -4664, -6519, 5246, 6048, 
---5789, -5531, 6283, 4968, -6728, -4368, 7118, 3730, -7452, -3065, 7725, 2374, -7938, -1666, 8086, 942, -8171, -214, 8189, -518, -8144, 1244, 8032, -1962, -7858, 2662, 7619, -3342, -7323, 3994, 
--6966, -4616, -6555, 5199, 6091, -5742, -5581, 6238, 5024, -6686, -4430, 7080, 3799, -7419, -3140, 7697, 2454, -7916, -1752, 8071, 1033, -8164, -309, 8190, -420, -8154, 1143, 8051, -1859, -7887, 
--2559, 7659, -3239, -7373, 3892, 7027, -4517, -6627, 5103, 6173, -5652, -5674, 6154, 5127, -6609, -4543, 7010, 3921, -7358, -3270, 7647, 2592, -7877, -1896, 8044, 1183, -8150, -464, 8190, -262, 
---8168, 983, 8080, -1698, -7931, 2397, 7718, -3080, -7447, 3737, 7116, -4366, -6732, 4959, 6293, -5515, -5808, 6027, 5275, -6493, -4704, 6907, 4094, -7268, -3454, 7572, 2786, -7818, -2099, 8002, 
--1393, -8126, -679, 8184, -43, -8182, 761, 8114, -1476, -7985, 2177, 7792, -2863, -7542, 3525, 7231, -4161, -6866, 4763, 6447, -5331, -5980, 5855, 5465, -6335, -4910, 6765, 4316, -7145, -3690, 
--7467, 3034, -7734, -2358, 7940, 1661, -8086, -953, 8169, 237, -8191, 479, 8148, -1194, -8044, 1896, 7877, -2587, -7652, 3255, 7366, -3900, -7026, 4513, 6631, -5094, -6187, 5633, 5694, -6132, 
---5159, 6581, 4584, -6982, -3975, 7328, 3335, -7620, -2671, 7852, 1985, -8026, -1286, 8137, 576, -8189, 136, 8176, -850, -8103, 1554, 7966, -2249, -7772, 2924, 7516, -3579, -7206, 4205, 6839, 
---4801, -6422, 5358, 5955, -5877, -5446, 6349, 4893, -6775, -4306, 7148, 3684, -7469, -3036, 7732, 2364, -7938, -1677, 8082, 974, -8168, -267, 8190, -444, -8153, 1149, 8052, -1848, -7893, 2531, 
--7673, -3196, -7397, 3836, 7064, -4448, -6680, 5025, 6244, -5566, -5764, 6064, 5238, -6518, -4676, 6921, 4077, -7274, -3450, 7571, 2795, -7813, -2121, 7995, 1430, -8120, -730, 8182, 23, -8185, 
--682, 8125, -1383, -8007, 2072, 7827, -2748, -7591, 3401, 7297, -4031, -6951, 4628, 6552, -5193, -6106, 5718, 5613, -6201, -5081, 6637, 4509, -7026, -3906, 7361, 3272, -7643, -2616, 7867, 1939, 
---8034, -1251, 8141, 551, -8189, 151, 8175, -854, -8103, 1548, 7969, -2232, -7779, 2898, 7529, -3544, -7227, 4163, 6869, -4752, -6463, 5304, 6008, -5820, -5511, 6290, 4971, -6717, -4398, 7092, 
--3790, -7417, -3157, 7686, 2499, -7901, -1825, 8055, 1135, -8153, -440, 8190, -260, -8169, 957, 8086, -1648, -7947, 2324, 7747, -2986, -7494, 3624, 7184, -4238, -6824, 4818, 6412, -5365, -5956, 
--5872, 5455, -6337, -4917, 6754, 4341, -7125, -3735, 7442, 3101, -7706, -2447, 7913, 1773, -8065, -1089, 8157, 395, -8191, 300, 8165, -994, -8081, 1679, 7938, -2354, -7739, 3010, 7483, -3645, 
---7175, 4253, 6813, -4831, -6405, 5373, 5948, -5878, -5452, 6339, 4914, -6756, -4343, 7122, 3739, -7440, -3110, 7702, 2458, -7911, -1790, 8061, 1107, -8156, -419, 8190, -274, -8168, 963, 8086, 
---1647, -7948, 2317, 7751, -2972, -7501, 3604, 7196, -4212, -6842, 4788, 6437, -5332, -5989, 5835, 5496, -6299, -4967, 6717, 4400, -7088, -3804, 7407, 3180, -7676, -2535, 7888, 1870, -8047, -1195, 
--8146, 509, -8190, 179, 8174, -867, -8102, 1546, 7971, -2217, -7786, 2869, 7544, -3503, -7251, 4111, 6905, -4691, -6513, 5236, 6073, -5746, -5592, 6214, 5070, -6640, -4515, 7017, 3927, -7347, 
---3312, 7623, 2673, -7848, -2018, 8016, 1346, -8129, -667, 8184, -18, -8184, 701, 8124, -1381, -8010, 2049, 7837, -2704, -7613, 3339, 7333, -3952, -7004, 4535, 6625, -5089, -6201, 5605, 5733, 
---6084, -5227, 6519, 4683, -6910, -4108, 7251, 3503, -7544, -2876, 7782, 2227, -7969, -1565, 8098, 891, -8173, -212, 8189, -470, -8151, 1146, 8055, -1816, -7905, 2472, 7699, -3112, -7442, 3729, 
--7131, -4322, -6773, 4883, 6367, -5412, -5920, 5902, 5429, -6353, -4904, 6758, 4343, -7119, -3754, 7429, 3138, -7690, -2502, 7896, 1847, -8050, -1182, 8147, 508, -8190, 169, 8175, -845, -8106, 
--1514, 7980, -2175, -7801, 2818, 7567, -3444, -7284, 4044, 6949, -4619, -6569, 5160, 6143, -5667, -5676, 6134, 5170, -6561, -4630, 6942, 4057, -7277, -3459, 7561, 2835, -7795, -2194, 7975, 1537, 
---8102, -871, 8173, 198, -8190, 474, 8150, -1145, -8057, 1806, 7908, -2457, -7707, 3089, 7452, -3702, -7149, 4288, 6797, -4846, -6400, 5370, 5958, -5860, -5479, 6308, 4961, -6716, -4412, 7076, 
--3831, -7391, -3227, 7654, 2599, -7868, -1956, 8027, 1298, -8134, -634, 8185, -37, -8183, 705, 8124, -1370, -8014, 2023, 7847, -2665, -7631, 3288, 7361, -3889, -7045, 4463, 6679, -5009, -6272, 
--5520, 5821, -5996, -5333, 6429, 4808, -6822, -4253, 7167, 3668, -7467, -3061, 7715, 2432, -7914, -1789, 8059, 1132, -8152, -470, 8189, -197, -8174, 860, 8103, -1520, -7981, 2167, 7804, -2802, 
---7578, 3416, 7299, -4009, -6975, 4574, 6603, -5111, -6189, 5612, 5733, -6078, -5242, 6501, 4714, -6884, -4157, 7220, 3571, -7510, -2964, 7749, 2336, -7939, -1695, 8075, 1041, -8161, -382, 8190, 
---281, -8169, 941, 8092, -1595, -7964, 2238, 7782, -2867, -7552, 3475, 7270, -4063, -6943, 4622, 6569, -5153, -6155, 5648, 5699, -6109, -5207, 6527, 4680, -6905, -4125, 7236, 3542, -7523, -2937, 
--7758, 2312, -7945, -1674, 8079, 1023, -8162, -368, 8190, -291, -8168, 947, 8091, -1598, -7964, 2236, 7783, -2862, -7554, 3467, 7275, -4052, -6951, 4608, 6581, -5137, -6170, 5631, 5718, -6090, 
---5231, 6508, 4708, -6886, -4158, 7218, 3579, -7505, -2980, 7743, 2359, -7932, -1726, 8069, 1080, -8157, -429, 8190, -227, -8173, 878, 8102, -1526, -7981, 2162, 7807, -2787, -7586, 3391, 7314, 
---3975, -6998, 4532, 6636, -5062, -6234, 5558, 5790, -6020, -5311, 6442, 4797, -6825, -4255, 7163, 3684, -7457, -3092, 7702, 2478, -7900, -1851, 8046, 1211, -8143, -565, 8187, -87, -8181, 735, 
--8122, -1381, -8013, 2016, 7852, -2640, -7644, 3245, 7385, -3832, -7083, 4392, 6733, -4927, -6344, 5428, 5913, -5898, -5447, 6328, 4945, -6720, -4414, 7069, 3854, -7375, -3272, 7632, 2668, -7844, 
---2049, 8005, 1415, -8118, -775, 8178, 128, -8189, 517, 8147, -1161, -8057, 1796, 7914, -2421, -7724, 3029, 7484, -3620, -7200, 4186, 6869, -4729, -6498, 5239, 6084, -5719, -5635, 6162, 5149, 
---6568, -4634, 6931, 4087, -7254, -3518, 7529, 2925, -7760, -2317, 7941, 1692, -8075, -1059, 8157, 418, -8191, 224, 8172, -866, -8105, 1501, 7987, -2128, -7821, 2740, 7605, -3337, -7345, 3911, 
--7037, -4463, -6689, 4986, 6298, -5480, -5870, 5938, 5405, -6362, -4908, 6744, 4380, -7088, -3827, 7386, 3249, -7641, -2653, 7847, 2040, -8007, -1416, 8116, 781, -8178, -144, 8189, -495, -8151, 
--1130, 8062, -1759, -7926, 2375, 7740, -2979, -7509, 3563, 7231, -4127, -6910, 4663, 6547, -5174, -6145, 5650, 5705, -6095, -5232, 6501, 4726, -6869, -4194, 7193, 3634, -7477, -3055, 7713, 2455, 
---7904, -1843, 8046, 1218, -8142, -587, 8186, -48, -8183, 681, 8130, -1312, -8029, 1933, 7878, -2544, -7682, 3137, 7439, -3714, -7152, 4266, 6822, -4794, -6452, 5292, 6042, -5760, -5598, 6191, 
--5119, -6588, -4611, 6942, 4074, -7258, -3515, 7528, 2934, -7755, -2337, 7935, 1724, -8068, -1103, 8152, 474, -8190, 156, 8177, -786, -8117, 1410, 8008, -2027, -7853, 2630, 7650, -3220, -7403, 
--3788, 7111, -4335, -6779, 4855, 6405, -5348, -5995, 5807, 5548, -6234, -5071, 6622, 4562, -6973, -4028, 7281, 3469, -7548, -2891, 7769, 2295, -7945, -1688, 8074, 1068, -8156, -445, 8189, -183, 
---8177, 807, 8114, -1429, -8006, 2040, 7849, -2641, -7648, 3224, 7400, -3790, -7112, 4332, 6780, -4851, -6411, 5339, 6003, -5798, -5562, 6221, 5086, -6610, -4583, 6958, 4052, -7268, -3499, 7533, 
--2925, -7757, -2335, 7934, 1730, -8067, -1118, 8151, 497, -8189, 125, 8179, -748, -8123, 1364, 8018, -1974, -7870, 2570, 7673, -3154, -7435, 3717, 7152, -4261, -6830, 4778, 6466, -5269, -6068, 
--5728, 5633, -6156, -5168, 6546, 4671, -6901, -4150, 7214, 3603, -7488, -3037, 7716, 2452, -7903, -1856, 8042, 1247, -8137, -633, 8184, 14, -8186, 603, 8140, -1219, -8049, 1825, 7910, -2423, 
---7728, 3005, 7501, -3571, -7232, 4115, 6921, -4638, -6573, 5132, 6185, -5599, -5765, 6032, 5310, -6432, -4827, 6794, 4315, -7120, -3781, 7403, 3223, -7646, -2650, 7844, 2059, -8000, -1460, 8109, 
--850, -8173, -237, 8190, -378, -8163, 989, 8088, -1597, -7969, 2193, 7804, -2779, -7597, 3347, 7345, -3898, -7054, 4425, 6722, -4929, -6354, 5403, 5949, -5849, -5513, 6260, 5044, -6638, -4549, 
--6977, 4027, -7279, -3484, 7538, 2921, -7757, -2343, 7930, 1750, -8062, -1150, 8147, 541, -8188, 68, 8182, -678, -8132, 1283, 8036, -1882, -7897, 2469, 7712, -3044, -7487, 3600, 7218, -4138, 
---6911, 4650, 6565, -5139, -6184, 5598, 5767, -6027, -5320, 6421, 4843, -6781, -4341, 7102, 3813, -7386, -3266, 7627, 2699, -7828, -2120, 7985, 1528, -8099, -929, 8166, 323, -8191, 282, 8170, 
---887, -8105, 1486, 7994, -2078, -7841, 2656, 7644, -3222, -7407, 3768, 7128, -4296, -6812, 4798, 6456, -5275, -6068, 5722, 5645, -6139, -5194, 6521, 4712, -6869, -4207, 7178, 3677, -7450, -3129, 
--7679, 2563, -7869, -1985, 8014, 1394, -8118, -798, 8175, 196, -8191, 405, 8160, -1005, -8087, 1598, 7969, -2184, -7810, 2757, 7606, -3316, -7364, 3855, 7080, -4375, -6760, 4870, 6403, -5340, 
---6012, 5779, 5588, -6189, -5136, 6564, 4654, -6906, -4150, 7209, 3622, -7475, -3076, 7698, 2512, -7883, -1937, 8024, 1350, -8123, -758, 8178, 160, -8190, 437, 8157, -1033, -8083, 1621, 7964, 
---2203, -7804, 2771, 7601, -3326, -7360, 3861, 7078, -4377, -6760, 4868, 6405, -5335, -6018, 5772, 5597, -6180, -5149, 6553, 4672, -6894, -4172, 7196, 3648, -7462, -3107, 7686, 2549, -7872, -1978, 
--8015, 1396, -8117, -809, 8174, 215, -8191, 378, 8163, -970, -8094, 1555, 7980, -2134, -7826, 2699, 7630, -3252, -7396, 3786, 7121, -4302, -6811, 4793, 6464, -5261, -6085, 5699, 5672, -6110, 
---5232, 6487, 4763, -6831, -4272, 7138, 3756, -7410, -3223, 7641, 2671, -7835, -2108, 7986, 1531, -8097, -949, 8164, 361, -8191, 227, 8174, -816, -8116, 1399, 8015, -1976, -7874, 2541, 7690, 
---3094, -7469, 3629, 7207, -4148, -6911, 4642, 6577, -5115, -6211, 5559, 5811, -5977, -5384, 6362, 4927, -6716, -4447, 7033, 3943, -7316, -3420, 7560, 2878, -7767, -2324, 7932, 1755, -8059, -1180, 
--8142, 598, -8186, -14, 8186, -572, -8146, 1152, 8063, -1728, -7940, 2294, 7776, -2849, -7574, 3388, 7331, -3912, -7054, 4413, 6738, -4894, -6391, 5348, 6009, -5776, -5599, 6174, 5159, -6542, 
---4695, 6874, 4205, -7174, -3697, 7436, 3167, -7662, -2624, 7847, 2066, -7995, -1500, 8100, 924, -8167, -346, 8190, -235, -8175, 814, 8116, -1389, -8019, 1956, 7879, -2515, -7702, 3059, 7485, 
---3590, -7232, 4100, 6941, -4592, -6617, 5058, 6259, -5502, -5871, 5915, 5453, -6301, -5009, 6654, 4538, -6975, -4047, 7259, 3534, -7509, -3006, 7720, 2461, -7895, -1906, 8028, 1340, -8123, -769, 
--8176, 192, -8191, 383, 8163, -958, -8097, 1526, 7988, -2088, -7843, 2638, 7656, -3177, -7434, 3698, 7174, -4202, -6880, 4684, 6550, -5144, -6191, 5577, 5799, -5985, -5380, 6361, 4934, -6707, 
---4465, 7019, 3973, -7298, -3463, 7539, 2935, -7745, -2394, 7912, 1840, -8041, -1279, 8130, 711, -8180, -140, 8189, -432, -8160, 1001, 8089, -1566, -7981, 2122, 7832, -2669, -7647, 3200, 7423, 
---3719, -7165, 4216, 6871, -4696, -6545, 5150, 6185, -5581, -5798, 5984, 5381, -6359, -4940, 6701, 4474, -7013, -3988, 7289, 3480, -7531, -2959, 7736, 2421, -7905, -1874, 8034, 1316, -8126, -754, 
--8177, 186, -8191, 380, 8164, -947, -8099, 1506, 7994, -2060, -7852, 2602, 7671, -3134, -7456, 3648, 7203, -4147, -6917, 4624, 6597, -5080, -6247, 5510, 5866, -5916, -5459, 6292, 5024, -6639, 
---4567, 6953, 4087, -7235, -3590, 7482, 3073, -7694, -2545, 7868, 2002, -8007, -1452, 8106, 894, -8168, -333, 8190, -231, -8176, 791, 8120, -1350, -8028, 1900, 7897, -2443, -7730, 2972, 7526, 
---3489, -7287, 3988, 7013, -4470, -6708, 4928, 6369, -5365, -6003, 5775, 5606, -6160, -5186, 6514, 4739, -6839, -4273, 7130, 3785, -7390, -3281, 7613, 2760, -7802, -2228, 7953, 1684, -8069, -1135, 
--8146, 578, -8186, -21, 8186, -538, -8151, 1092, 8075, -1643, -7964, 2185, 7815, -2718, -7631, 3236, 7410, -3741, -7156, 4226, 6868, -4694, -6550, 5138, 6200, -5560, -5823, 5955, 5418, -6323, 
---4990, 6661, 4537, -6970, -4066, 7244, 3574, -7487, -3067, 7694, 2545, -7868, -2013, 8003, 1471, -8103, -923, 8165, 370, -8191, 183, 8178, -736, -8129, 1285, 8041, -1829, -7919, 2362, 7758, 
---2887, -7564, 3396, 7334, -3892, -7073, 4368, 6777, -4826, -6453, 5260, 6098, -5671, -5717, 6055, 5308, -6413, -4878, 6741, 4423, -7039, -3951, 7304, 3459, -7537, -2953, 7735, 2433, -7899, -1903, 
--8026, 1364, -8118, -820, 8172, 271, -8191, 277, 8172, -826, -8118, 1369, 8025, -1908, -7898, 2435, 7734, -2954, -7537, 3457, 7305, -3947, -7042, 4417, 6746, -4869, -6422, 5297, 6067, -5703, 
---5687, 6081, 5280, -6435, -4852, 6758, 4400, -7052, -3931, 7313, 3442, -7543, -2941, 7738, 2424, -7901, -1899, 8026, 1364, -8118, -825, 8172, 280, -8191, 263, 8173, -808, -8120, 1346, 8030, 
---1880, -7906, 2404, 7745, -2919, -7553, 3419, 7325, -3906, -7067, 4374, 6776, -4824, -6458, 5250, 6109, -5656, -5735, 6035, 5335, -6389, -4913, 6713, 4468, -7009, -4006, 7273, 3524, -7507, -3029, 
--7706, 2519, -7873, -2001, 8004, 1471, -8102, -938, 8163, 398, -8190, 140, 8180, -680, -8136, 1215, 8055, -1747, -7941, 2269, 7791, -2782, -7609, 3282, 7392, -3769, -7145, 4237, 6866, -4690, 
---6559, 5119, 6222, -5529, -5860, 5912, 5471, -6272, -5060, 6603, 4626, -6908, -4175, 7180, 3703, -7424, -3218, 7633, 2717, -7812, -2207, 7956, 1685, -8067, -1159, 8142, 625, -8184, -91, 8189, 
---445, -8161, 977, 8096, -1506, -7999, 2027, 7865, -2541, -7701, 3042, 7501, -3532, -7272, 4005, 7010, -4463, -6720, 4899, 6400, -5317, -6055, 5710, 5683, -6081, -5288, 6424, 4870, -6741, -4433, 
--7028, 3975, -7287, -3503, 7514, 3014, -7710, -2515, 7872, 2003, -8003, -1486, 8099, 960, -8162, -432, 8189, -100, -8183, 628, 8142, -1156, -8068, 1677, 7958, -2193, -7818, 2697, 7642, -3192, 
---7437, 3672, 7199, -4138, -6933, 4584, 6636, -5013, -6313, 5419, 5963, -5805, -5590, 6164, 5192, -6500, -4774, 6806, 4335, -7086, -3879, 7335, 3406, -7555, -2922, 7742, 2423, -7899, -1916, 8021, 
--1400, -8112, -880, 8167, 354, -8191, 170, 8179, -696, -8135, 1217, 8056, -1734, -7946, 2242, 7802, -2743, -7627, 3231, 7419, -3706, -7183, 4165, 6915, -4608, -6622, 5031, 6299, -5434, -5953, 
--5814, 5580, -6171, -5187, 6501, 4771, -6807, -4338, 7082, 3885, -7331, -3419, 7548, 2937, -7736, -2445, 7891, 1942, -8016, -1432, 8106, 915, -8165, -397, 8189, -125, -8182, 644, 8141, -1162, 
---8068, 1673, 7960, -2180, -7823, 2675, 7652, -3162, -7453, 3634, 7221, -4092, -6963, 4533, 6675, -4956, -6362, 5358, 6022, -5741, -5659, 6098, 5273, -6432, -4867, 6739, 4440, -7020, -3997, 7272, 
--3537, -7496, -3064, 7689, 2578, -7853, -2084, 7983, 1579, -8084, -1071, 8150, 556, -8186, -41, 8188, -475, -8159, 988, 8096, -1498, -8002, 2001, 7875, -2497, -7719, 2981, 7531, -3455, -7315, 
--3914, 7068, -4359, -6796, 4784, 6494, -5193, -6170, 5578, 5819, -5944, -5447, 6285, 5053, -6602, -4640, 6892, 4208, -7156, -3761, 7390, 3298, -7598, -2824, 7773, 2337, -7920, -1843, 8034, 1340, 
---8119, -834, 8170, 323, -8191, 187, 8179, -698, -8136, 1204, 8060, -1707, -7955, 2202, 7817, -2689, -7650, 3164, 7452, -3629, -7227, 4078, 6973, -4512, -6693, 4927, 6386, -5325, -6057, 5700, 
--5702, -6055, -5327, 6384, 4930, -6691, -4516, 6970, 4083, -7224, -3636, 7448, 3174, -7646, -2701, 7812, 2217, -7950, -1726, 8056, 1227, -8133, -725, 8177, 219, -8191, 286, 8173, -792, -8125, 
--1292, 8044, -1790, -7935, 2278, 7793, -2760, -7624, 3229, 7424, -3687, -7198, 4129, 6943, -4558, -6663, 4967, 6357, -5359, -6028, 5728, 5675, -6078, -5303, 6403, 4908, -6705, -4498, 6980, 4068, 
---7231, -3626, 7452, 3168, -7648, -2700, 7812, 2220, -7949, -1734, 8054, 1240, -8131, -743, 8176, 242, -8191, 258, 8175, -759, -8129, 1254, 8052, -1747, -7946, 2232, 7809, -2709, -7644, 3175, 
--7450, -3630, -7229, 4070, 6980, -4496, -6707, 4904, 6408, -5295, -6086, 5664, 5741, -6015, -5376, 6341, 4989, -6645, -4586, 6923, 4165, -7177, -3730, 7402, 3279, -7602, -2819, 7772, 2346, -7916, 
---1867, 8028, 1380, -8113, -889, 8165, 393, -8190, 101, 8183, -598, -8148, 1090, 8081, -1579, -7987, 2061, 7861, -2537, -7709, 3002, 7526, -3457, -7319, 3898, 7082, -4326, -6823, 4737, 6536, 
---5132, -6228, 5506, 5895, -5862, -5543, 6195, 5169, -6507, -4779, 6793, 4369, -7057, -3946, 7293, 3506, -7505, -3056, 7687, 2594, -7844, -2124, 7971, 1645, -8070, -1162, 8139, 673, -8180, -183, 
--8190, -308, -8173, 797, 8124, -1284, -8048, 1765, 7942, -2241, -7809, 2707, 7646, -3165, -7458, 3609, 7241, -4042, -7001, 4459, 6734, -4862, -6445, 5246, 6131, -5612, -5797, 5957, 5441, -6282, 
---5068, 6583, 4675, -6862, -4268, 7115, 3844, -7344, -3408, 7546, 2959, -7723, -2501, 7870, 2032, -7992, -1559, 8084, 1078, -8149, -596, 8183, 109, -8190, 375, 8167, -860, -8117, 1340, 8037, 
---1816, -7930, 2285, 7794, -2747, -7633, 3197, 7443, -3638, -7229, 4064, 6988, -4478, -6724, 4874, 6436, -5254, -6127, 5615, 5795, -5957, -5445, 6277, 5074, -6577, -4687, 6852, 4283, -7105, -3866, 
--7332, 3433, -7535, -2991, 7710, 2537, -7860, -2076, 7981, 1607, -8076, -1134, 8142, 655, -8181, -176, 8190, -305, -8173, 783, 8126, -1260, -8054, 1731, 7951, -2197, -7824, 2654, 7667, -3104, 
---7487, 3540, 7279, -3967, -7048, 4378, 6791, -4775, -6514, 5154, 6212, -5518, -5891, 5860, 5548, -6185, -5189, 6486, 4810, -6767, -4417, 7024, 4007, -7258, -3586, 7465, 3150, -7650, -2707, 7806, 
--2252, -7938, -1792, 8041, 1324, -8119, -854, 8167, 379, -8190, 95, 8184, -571, -8152, 1042, 8090, -1512, -8004, 1974, 7888, -2432, -7749, 2879, 7581, -3318, -7390, 3744, 7173, -4160, -6934, 
--4559, 6669, -4945, -6385, 5313, 6077, -5665, -5752, 5995, 5405, -6308, -5043, 6597, 4662, -6867, -4267, 7111, 3857, -7334, -3436, 7531, 3002, -7704, -2560, 7851, 2108, -7973, -1651, 8067, 1187, 
---8136, -721, 8176, 251, -8191, 217, 8178, -687, -8140, 1152, 8073, -1616, -7981, 2071, 7862, -2522, -7718, 2963, 7548, -3395, -7355, 3814, 7136, -4223, -6896, 4616, 6631, -4995, -6347, 5356, 
--6041, -5702, -5717, 6027, 5372, -6334, -5013, 6618, 4635, -6883, -4244, 7123, 3838, -7343, -3421, 7536, 2992, -7707, -2555, 7851, 2108, -7972, -1656, 8065, 1198, -8134, -737, 8175, 273, -8191, 
--190, 8180, -655, -8144, 1115, 8079, -1573, -7991, 2024, 7876, -2471, -7737, 2907, 7572, -3336, -7384, 3752, 7171, -4158, -6938, 4548, 6680, -4926, -6403, 5286, 6104, -5631, -5788, 5957, 5451, 
---6265, -5100, 6551, 4730, -6818, -4348, 7061, 3950, -7284, -3541, 7482, 3120, -7659, -2691, 7809, 2251, -7936, -1807, 8036, 1355, -8113, -902, 8163, 443, -8189, 14, 8187, -474, -8161, 930, 
--8108, -1384, -8032, 1832, 7928, -2276, -7802, 2711, 7650, -3140, -7476, 3556, 7276, -3963, -7056, 4355, 6812, -4736, -6549, 5100, 6264, -5450, -5962, 5781, 5639, -6096, -5301, 6390, 4944, -6665, 
---4575, 6919, 4189, -7153, -3793, 7362, 3383, -7551, -2965, 7714, 2536, -7856, -2102, 7972, 1659, -8065, -1213, 8131, 762, -8174, -310, 8190, -144, -8183, 595, 8149, -1047, -8092, 1493, 8009, 
---1936, -7903, 2372, 7771, -2801, -7618, 3221, 7439, -3632, -7240, 4030, 7017, -4417, -6774, 4789, 6510, -5149, -6228, 5490, 5925, -5817, -5606, 6124, 5268, -6414, -4917, 6683, 4549, -6934, -4169, 
--7162, 3775, -7370, -3372, 7554, 2957, -7717, -2535, 7855, 2104, -7971, -1669, 8061, 1227, -8130, -783, 8171, 336, -8191, 111, 8184, -559, -8154, 1003, 8098, -1446, -8021, 1882, 7917, -2315, 
---7792, 2739, 7641, -3156, -7471, 3562, 7276, -3959, -7061, 4342, 6824, -4714, -6569, 5070, 6292, -5413, -5999, 5738, 5687, -6047, -5360, 6337, 5015, -6610, -4657, 6862, 4285, -7095, -3901, 7305, 
--3505, -7496, -3100, 7662, 2684, -7809, -2263, 7930, 1834, -8030, -1401, 8105, 962, -8158, -523, 8185, 80, -8190, 361, 8170, -802, -8128, 1239, 8060, -1674, -7971, 2102, 7857, -2526, -7722, 
--2940, 7563, -3348, -7384, 3744, 7181, -4131, -6961, 4503, 6718, -4865, -6458, 5210, 6177, -5542, -5881, 5857, 5566, -6156, -5238, 6435, 4892, -6698, -4535, 6940, 4163, -7163, -3781, 7364, 3386, 
---7546, -2984, 7705, 2572, -7843, -2154, 7957, 1729, -8050, -1300, 8118, 867, -8166, -433, 8188, -4, -8188, 439, 8164, -874, -8119, 1305, 8048, -1734, -7957, 2156, 7842, -2573, -7706, 2981, 
--7547, -3382, -7368, 3772, 7167, -4153, -6948, 4520, 6708, -4876, -6451, 5217, 6174, -5545, -5881, 5855, 5571, -6150, -5247, 6426, 4906, -6686, -4554, 6926, 4188, -7148, -3812, 7348, 3423, -7529, 
---3027, 7688, 2621, -7827, -2210, 7942, 1791, -8038, -1369, 8109, 942, -8159, -514, 8185, 83, -8190, 346, 8171, -776, -8132, 1201, 8068, -1626, -7983, 2043, 7875, -2457, -7748, 2861, 7597, 
---3260, -7427, 3648, 7235, -4027, -7026, 4393, 6795, -4749, -6548, 5090, 6281, -5419, -6000, 5731, 5700, -6029, -5386, 6309, 5056, -6574, -4715, 6818, 4359, -7046, -3993, 7253, 3615, -7442, -3229, 
--7609, 2833, -7757, -2431, 7882, 2020, -7988, -1607, 8070, 1187, -8133, -766, 8172, 342, -8190, 81, 8185, -506, -8160, 928, 8111, -1348, -8042, 1763, 7950, -2175, -7839, 2579, 7705, -2978, 
---7552, 3366, 7377, -3748, -7185, 4117, 6972, -4478, -6742, 4824, 6492, -5159, -6228, 5479, 5945, -5786, -5648, 6075, 5335, -6350, -5010, 6607, 4669, -6848, -4319, 7068, 3955, -7272, -3583, 7455, 
--3200, -7620, -2811, 7763, 2412, -7887, -2009, 7989, 1600, -8072, -1188, 8132, 771, -8172, -355, 8189, -65, -8187, 482, 8161, -899, -8117, 1312, 8049, -1723, -7962, 2128, 7852, -2529, -7725, 
--2921, 7575, -3307, -7408, 3683, 7220, -4051, -7015, 4406, 6790, -4752, -6550, 5084, 6291, -5404, -6018, 5708, 5727, -5999, -5424, 6273, 5105, -6532, -4776, 6773, 4432, -6998, -4079, 7204, 3714, 
---7392, -3341, 7560, 2959, -7711, -2570, 7839, 2174, -7950, -1774, 8038, 1368, -8108, -960, 8156, 548, -8184, -137, 8190, -276, -8177, 686, 8142, -1096, -8088, 1501, 8011, -1905, -7917, 2301, 
--7800, -2693, -7666, 3077, 7511, -3454, -7339, 3821, 7147, -4180, -6938, 4526, 6711, -4863, -6469, 5185, 6208, -5496, -5935, 5792, 5645, -6075, -5342, 6340, 5025, -6592, -4697, 6825, 4356, -7043, 
---4006, 7242, 3645, -7424, -3276, 7586, 2898, -7731, -2514, 7855, 2123, -7962, -1728, 8047, 1328, -8114, -926, 8158, 521, -8185, -116, 8190, -291, -8177, 695, 8141, -1099, -8088, 1498, 8013, 
---1896, -7920, 2286, 7806, -2673, -7675, 3051, 7523, -3423, -7355, 3785, 7168, -4140, -6965, 4482, 6743, -4815, -6507, 5134, 6253, -5443, -5986, 5737, 5703, -6018, -5408, 6283, 5098, -6534, -4778, 
--6768, 4445, -6987, -4103, 7187, 3750, -7372, -3390, 7537, 3019, -7686, -2644, 7815, 2261, -7926, -1874, 8017, 1481, -8090, -1087, 8142, 688, -8177, -290, 8190, -111, -8186, 509, 8160, -908, 
---8117, 1303, 8052, -1696, -7971, 2083, 7868, -2466, -7749, 2842, 7610, -3213, -7455, 3574, 7280, -3929, -7091, 4272, 6882, -4607, -6660, 4929, 6420, -5241, -6167, 5539, 5898, -5825, -5617, 6096, 
--5321, -6354, -5015, 6596, 4695, -6823, -4366, 7033, 4026, -7229, -3678, 7405, 3320, -7566, -2956, 7708, 2584, -7833, -2208, 7938, 1824, -8027, -1439, 8095, 1049, -8147, -658, 8177, 265, -8191, 
--128, 8184, -522, -8160, 912, 8115, -1302, -8054, 1687, 7972, -2070, -7874, 2446, 7756, -2818, -7622, 3181, 7469, -3539, -7301, 3887, 7114, -4228, -6913, 4557, 6695, -4877, -6463, 5184, 6215, 
---5482, -5955, 5764, 5680, -6036, -5393, 6291, 5093, -6534, -4783, 6761, 4461, -6974, -4131, 7169, 3790, -7350, -3442, 7512, 3085, -7659, -2723, 7787, 2353, -7900, -1980, 7992, 1600, -8069, -1220, 
--8126, 834, -8166, -449, 8187, 62, -8190, 324, 8174, -711, -8142, 1094, 8089, -1476, -8021, 1853, 7932, -2227, -7828, 2595, 7705, -2958, -7567, 3313, 7410, -3662, -7239, 4001, 7051, -4333, 
---6848, 4654, 6629, -4965, -6397, 5264, 6149, -5553, -5890, 5828, 5616, -6092, -5332, 6340, 5035, -6577, -4729, 6797, 4410, -7004, -4084, 7193, 3747, -7369, -3405, 7527, 3053, -7670, -2696, 7795, 
--2332, -7904, -1965, 7995, 1592, -8070, -1218, 8126, 839, -8166, -461, 8186, 80, -8191, 299, 8176, -679, -8145, 1056, 8095, -1432, -8030, 1803, 7946, -2171, -7846, 2533, 7728, -2892, -7595, 
--3242, 7445, -3587, -7280, 3922, 7098, -4250, -6903, 4567, 6691, -4877, -6468, 5174, 6228, -5462, -5978, 5736, 5713, -5999, -5438, 6248, 5150, -6486, -4853, 6708, 4544, -6918, -4228, 7110, 3901, 
---7290, -3568, 7453, 3225, -7602, -2878, 7732, 2523, -7849, -2165, 7947, 1801, -8030, -1435, 8095, 1064, -8144, -693, 8175, 319, -8190, 53, 8187, -427, -8169, 798, 8131, -1169, -8079, 1536, 
--8008, -1901, -7923, 2260, 7819, -2616, -7701, 2965, 7566, -3309, -7416, 3645, 7250, -3975, -7071, 4294, 6875, -4606, -6668, 4907, 6445, -5200, -6211, 5479, 5962, -5750, -5703, 6006, 5431, -6253, 
---5150, 6484, 4857, -6704, -4555, 6908, 4243, -7100, -3924, 7276, 3596, -7439, -3262, 7585, 2920, -7717, -2574, 7831, 2222, -7932, -1867, 8015, 1506, -8084, -1145, 8134, 779, -8170, -414, 8187, 
--47, -8190, 319, 8175, -685, -8145, 1048, 8098, -1411, -8036, 1769, 7956, -2125, -7862, 2475, 7750, -2821, -7626, 3160, 7484, -3494, -7330, 3819, 7159, -4139, -6976, 4448, 6777, -4750, -6567, 
--5040, 6342, -5323, -6107, 5593, 5858, -5854, -5599, 6101, 5328, -6338, -5049, 6560, 4757, -6772, -4459, 6968, 4150, -7152, -3835, 7320, 3511, -7476, -3182, 7616, 2845, -7742, -2505, 7852, 2158, 
---7948, -1809, 8026, 1454, -8091, -1099, 8139, 741, -8172, -383, 8188, 22, -8190, 336, 8174, -696, -8145, 1052, 8098, -1408, -8037, 1759, 7959, -2108, -7868, 2451, 7759, -2792, -7638, 3124, 
--7501, -3453, -7351, 3773, 7186, -4087, -7008, 4392, 6816, -4690, -6613, 4977, 6395, -5256, -6167, 5524, 5926, -5782, -5676, 6028, 5413, -6264, -5142, 6486, 4859, -6698, -4570, 6895, 4270, -7081, 
---3964, 7252, 3649, -7411, -3329, 7554, 3002, -7685, -2670, 7799, 2332, -7901, -1992, 7986, 1647, -8058, -1300, 8113, 949, -8155, -599, 8180, 246, -8191, 106, 8186, -459, -8167, 809, 8131, 
---1159, -8082, 1505, 8017, -1850, -7938, 2190, 7843, -2527, -7736, 2857, 7613, -3184, -7477, 3503, 7327, -3818, -7164, 4123, 6987, -4423, -6799, 4712, 6597, -4994, -6385, 5266, 6159, -5529, -5925, 
--5781, 5678, -6024, -5422, 6253, 5155, -6474, -4881, 6680, 4596, -6876, -4305, 7058, 4005, -7229, -3699, 7385, 3385, -7529, -3067, 7658, 2741, -7775, -2413, 7876, 2079, -7965, -1743, 8038, 1403, 
---8098, -1062, 8142, 717, -8173, -373, 8188, 27, -8190, 317, 8176, -662, -8149, 1004, 8106, -1346, -8050, 1684, 7978, -2020, -7895, 2350, 7795, -2678, -7684, 3000, 7557, -3317, -7419, 3627, 
--7266, -3932, -7102, 4229, 6924, -4519, -6736, 4800, 6535, -5074, -6324, 5337, 6100, -5592, -5868, 5836, 5624, -6071, -5372, 6294, 5109, -6508, -4839, 6708, 4559, -6899, -4273, 7075, 3978, -7241, 
---3678, 7393, 3371, -7534, -3059, 7660, 2741, -7774, -2420, 7874, 2093, -7961, -1764, 8033, 1431, -8093, -1098, 8138, 761, -8170, -424, 8187, 86, -8191, 251, 8180, -589, -8156, 924, 8117, 
---1259, -8067, 1590, 8000, -1920, -7922, 2244, 7829, -2567, -7725, 2883, 7605, -3196, -7475, 3501, 7331, -3803, -7176, 4095, 7008, -4383, -6829, 4662, 6638, -4934, -6437, 5196, 6224, -5451, -6002, 
--5695, 5769, -5931, -5528, 6155, 5277, -6371, -5018, 6574, 4750, -6769, -4476, 6950, 4192, -7121, -3904, 7278, 3607, -7426, -3307, 7559, 3000, -7682, -2689, 7789, 2373, -7887, -2055, 7969, 1731, 
---8040, -1407, 8096, 1079, -8140, -752, 8169, 421, -8187, -92, 8190, -239, -8182, 568, 8158, -897, -8123, 1223, 8072, -1549, -8011, 1870, 7935, -2189, -7848, 2503, 7747, -2815, -7635, 3120, 
--7509, -3422, -7373, 3716, 7223, -4006, -7064, 4288, 6891, -4564, -6710, 4831, 6516, -5092, -6314, 5343, 6100, -5587, -5878, 5821, 5645, -6046, -5405, 6261, 5155, -6467, -4899, 6660, 4633, -6845, 
---4363, 7018, 4083, -7181, -3799, 7330, 3508, -7470, -3213, 7597, 2911, -7713, -2607, 7815, 2296, -7907, -1985, 7984, 1669, -8051, -1352, 8103, 1031, -8145, -711, 8172, 388, -8188, -67, 8190, 
---257, -8181, 578, 8157, -899, -8123, 1217, 8074, -1535, -8015, 1849, 7941, -2161, -7858, 2468, 7760, -2773, -7652, 3071, 7531, -3367, -7400, 3655, 7257, -3940, -7104, 4216, 6938, -4488, -6764, 
--4751, 6578, -5008, -6384, 5256, 6178, -5497, -5965, 5728, 5742, -5952, -5511, 6165, 5271, -6371, -5025, 6565, 4769, -6751, -4508, 6925, 4239, -7090, -3965, 7242, 3684, -7386, -3400, 7516, 3108, 
---7637, -2814, 7745, 2514, -7843, -2213, 7927, 1906, -8002, -1599, 8062, 1287, -8113, -976, 8149, 662, -8176, -349, 8188, 33, -8191, 280, 8179, -595, -8157, 907, 8121, -1219, -8076, 1527, 
--8016, -1835, -7947, 2137, 7864, -2439, -7772, 2735, 7667, -3028, -7552, 3315, 7425, -3599, -7289, 3876, 7140, -4149, -6983, 4413, 6814, -4674, -6638, 4925, 6450, -5171, -6254, 5407, 6048, -5637, 
---5835, 5858, 5613, -6071, -5384, 6274, 5145, -6470, -4902, 6654, 4649, -6830, -4392, 6995, 4127, -7152, -3858, 7297, 3582, -7433, -3303, 7556, 3018, -7671, -2730, 7772, 2437, -7865, -2143, 7944, 
--1843, -8014, -1544, 8071, 1240, -8119, -937, 8153, 630, -8178, -325, 8189, 18, -8190, 287, 8179, -594, -8157, 898, 8123, -1202, -8079, 1502, 8022, -1802, -7956, 2097, 7877, -2391, -7789, 
--2680, 7688, -2967, -7579, 3247, 7458, -3525, -7328, 3796, 7186, -4063, -7037, 4323, 6875, -4578, -6707, 4825, 6527, -5068, -6341, 5301, 6144, -5529, -5941, 5747, 5728, -5960, -5510, 6162, 5282, 
---6357, -5049, 6542, 4807, -6720, -4561, 6886, 4307, -7046, -4049, 7193, 3784, -7333, -3516, 7461, 3242, -7581, -2965, 7688, 2683, -7787, -2399, 7874, 2110, -7952, -1821, 8018, 1527, -8074, -1233, 
--8118, 936, -8153, -640, 8176, 342, -8189, -45, 8190, -254, -8182, 550, 8161, -848, -8131, 1142, 8088, -1436, -8037, 1726, 7974, -2016, -7902, 2301, 7818, -2585, -7725, 2863, 7621, -3139, 
---7508, 3409, 7384, -3677, -7253, 3937, 7110, -4194, -6960, 4444, 6799, -4689, -6631, 4927, 6453, -5160, -6269, 5384, 6075, -5603, -5875, 5812, 5665, -6016, -5451, 6211, 5228, -6399, -5000, 6576, 
--4764, -6748, -4524, 6908, 4276, -7062, -4025, 7204, 3767, -7340, -3507, 7463, 3240, -7580, -2971, 7684, 2697, -7781, -2422, 7866, 2141, -7943, -1860, 8008, 1575, -8065, -1291, 8110, 1003, -8146, 
---715, 8171, 425, -8187, -137, 8190, -153, -8186, 441, 8170, -730, -8145, 1016, 8108, -1303, -8063, 1585, 8006, -1868, -7942, 2146, 7865, -2423, -7781, 2696, 7686, -2966, -7583, 3231, 7468, 
---3493, -7347, 3750, 7215, -4003, -7076, 4249, 6926, -4492, -6771, 4728, 6605, -4959, -6433, 5182, 6251, -5401, -6064, 5611, 5868, -5816, -5667, 6012, 5457, -6203, -5242, 6384, 5020, -6559, -4793, 
--6724, 4559, -6883, -4322, 7031, 4078, -7173, -3831, 7305, 3577, -7429, -3322, 7543, 3060, -7650, -2798, 7745, 2530, -7833, -2261, 7910, 1988, -7980, -1714, 8037, 1437, -8088, -1161, 8127, 881, 
---8158, -602, 8177, 321, -8190, -41, 8190, -240, -8183, 519, 8164, -799, -8138, 1076, 8100, -1353, -8055, 1627, 7998, -1900, -7935, 2169, 7860, -2438, -7778, 2701, 7685, -2963, -7585, 3220, 
--7475, -3475, -7358, 3723, 7231, -3969, -7098, 4208, 6954, -4445, -6805, 4674, 6646, -4899, -6481, 5117, 6308, -5331, -6129, 5537, 5941, -5738, -5749, 5930, 5548, -6118, -5344, 6297, 5131, -6470, 
---4915, 6634, 4691, -6792, -4464, 6941, 4231, -7084, -3995, 7216, 3752, -7343, -3508, 7459, 3257, -7569, -3006, 7668, 2749, -7761, -2491, 7843, 2229, -7918, -1966, 7983, 1700, -8040, -1433, 8087, 
--1164, -8127, -895, 8155, 623, -8177, -353, 8188, 81, -8191, 189, 8184, -461, -8170, 730, 8145, -1000, -8113, 1267, 8070, -1534, -8020, 1797, 7960, -2060, -7893, 2319, 7816, -2577, -7732, 
--2830, 7638, -3082, -7538, 3328, 7428, -3573, -7312, 3811, 7186, -4048, -7055, 4277, 6914, -4504, -6768, 4724, 6612, -4941, -6452, 5151, 6283, -5357, -6110, 5555, 5928, -5748, -5742, 5934, 5548, 
---6116, -5350, 6288, 5145, -6456, -4937, 6615, 4721, -6769, -4503, 6914, 4278, -7053, -4051, 7183, 3818, -7308, -3583, 7422, 3342, -7531, -3100, 7630, 2854, -7723, -2606, 7806, 2354, -7883, -2101, 
--7949, 1845, -8010, -1589, 8059, 1329, -8103, -1071, 8136, 809, -8163, -549, 8180, 286, -8190, -25, 8190, -237, -8183, 497, 8166, -759, -8143, 1017, 8110, -1276, -8070, 1532, 8020, -1788, 
---7965, 2040, 7899, -2292, -7827, 2539, 7746, -2786, -7658, 3027, 7562, -3267, -7459, 3502, 7348, -3735, -7231, 3963, 7104, -4188, -6973, 4407, 6834, -4623, -6689, 4832, 6536, -5039, -6379, 5238, 
--6213, -5435, -6043, 5623, 5866, -5808, -5685, 5985, 5496, -6158, -5305, 6323, 5106, -6484, -4904, 6636, 4696, -6784, -4486, 6923, 4269, -7057, -4050, 7182, 3825, -7302, -3599, 7413, 3368, -7518, 
---3135, 7615, 2898, -7706, -2660, 7787, 2418, -7863, -2175, 7929, 1929, -7990, -1683, 8041, 1434, -8086, -1185, 8122, 934, -8151, -684, 8172, 431, -8186, -180, 8190, -73, -8189, 323, 8178, 
---575, -8162, 825, 8135, -1075, -8103, 1322, 8062, -1570, -8015, 1814, 7958, -2058, -7897, 2298, 7825, -2538, -7749, 2773, 7664, -3007, -7573, 3237, 7474, -3465, -7369, 3688, 7256, -3909, -7139, 
--4125, 7013, -4338, -6882, 4546, 6744, -4751, -6601, 4949, 6450, -5145, -6296, 5334, 6134, -5520, -5968, 5699, 5796, -5875, -5620, 6043, 5437, -6207, -5252, 6364, 5059, -6517, -4865, 6662, 4664, 
---6803, -4461, 6935, 4253, -7064, -4042, 7183, 3827, -7299, -3610, 7406, 3388, -7508, -3165, 7601, 2937, -7689, -2710, 7769, 2477, -7844, -2245, 7909, 2009, -7970, -1774, 8022, 1535, -8068, -1297, 
--8106, 1056, -8138, -817, 8161, 574, -8179, -334, 8188, 91, -8191, 149, 8186, -391, -8176, 631, 8156, -872, -8131, 1110, 8098, -1348, -8059, 1584, 8012, -1820, -7959, 2052, 7898, -2284, 
---7833, 2512, 7758, -2740, -7679, 2963, 7592, -3185, -7500, 3403, 7400, -3619, -7295, 3831, 7183, -4040, -7067, 4245, 6942, -4447, -6814, 4644, 6679, -4838, -6540, 5027, 6393, -5212, -6243, 5392, 
--6087, -5569, -5927, 5739, 5760, -5906, -5591, 6066, 5415, -6223, -5237, 6372, 5053, -6518, -4867, 6657, 4675, -6792, -4481, 6920, 4282, -7043, -4081, 7159, 3876, -7271, -3669, 7375, 3457, -7474, 
---3245, 7566, 3028, -7653, -2811, 7732, 2590, -7807, -2369, 7873, 2145, -7935, -1920, 7989, 1693, -8038, -1466, 8078, 1236, -8114, -1008, 8142, 777, -8165, -547, 8179, 315, -8189, -85, 8190, 
---146, -8187, 376, 8176, -607, -8160, 835, 8135, -1064, -8106, 1291, 8069, -1518, -8028, 1741, 7978, -1966, -7924, 2186, 7862, -2407, -7796, 2623, 7722, -2840, -7643, 3051, 7557, -3263, -7468, 
--3469, 7370, -3675, -7269, 3876, 7161, -4076, -7049, 4270, 6929, -4463, -6807, 4650, 6677, -4836, -6545, 5015, 6405, -5193, -6263, 5365, 6114, -5534, -5963, 5697, 5805, -5858, -5645, 6012, 5479, 
---6163, -5311, 6308, 5137, -6450, -4961, 6585, 4780, -6716, -4598, 6841, 4410, -6962, -4221, 7076, 4027, -7187, -3832, 7291, 3633, -7390, -3433, 7483, 3228, -7571, -3024, 7652, 2815, -7730, -2607, 
--7799, 2395, -7865, -2183, 7923, 1968, -7977, -1753, 8024, 1536, -8066, -1320, 8101, 1100, -8131, -883, 8154, 662, -8173, -444, 8184, 223, -8191, -5, 8190, -216, -8185, 434, 8172, -653, 
---8156, 870, 8132, -1088, -8104, 1303, 8068, -1519, -8029, 1732, 7981, -1945, -7931, 2155, 7873, -2365, -7811, 2571, 7742, -2777, -7669, 2979, 7589, -3181, -7506, 3378, 7416, -3575, -7323, 3767, 
--7222, -3958, -7119, 4145, 7009, -4330, -6896, 4510, 6777, -4689, -6655, 4863, 6526, -5035, -6395, 5201, 6258, -5366, -6119, 5525, 5973, -5682, -5826, 5833, 5673, -5982, -5518, 6124, 5358, -6265, 
---5196, 6399, 5029, -6531, -4860, 6656, 4687, -6778, -4512, 6894, 4333, -7007, -4152, 7113, 3968, -7217, -3782, 7313, 3593, -7407, -3403, 7494, 3209, -7577, -3015, 7654, 2818, -7727, -2620, 7793, 
--2419, -7856, -2219, 7912, 2016, -7965, -1813, 8010, 1607, -8052, -1403, 8087, 1196, -8118, -990, 8142, 782, -8163, -575, 8177, 366, -8187, -160, 8190, -49, -8190, 255, 8183, -464, -8172, 
--669, 8154, -876, -8133, 1080, 8105, -1286, -8073, 1488, 8035, -1691, -7993, 1891, 7945, -2092, -7893, 2289, 7835, -2486, -7774, 2680, 7705, -2873, -7635, 3063, 7557, -3253, -7477, 3438, 7390, 
---3624, -7301, 3804, 7205, -3985, -7107, 4160, 7003, -4335, -6896, 4505, 6784, -4674, -6669, 4838, 6548, -5001, -6426, 5159, 6297, -5315, -6167, 5466, 6031, -5616, -5894, 5760, 5751, -5902, -5607, 
--6039, 5458, -6174, -5308, 6303, 5152, -6430, -4996, 6551, 4835, -6671, -4673, 6784, 4506, -6895, -4339, 6999, 4168, -7102, -3996, 7198, 3820, -7292, -3644, 7379, 3464, -7464, -3284, 7543, 3100, 
---7619, -2917, 7688, 2730, -7755, -2544, 7816, 2355, -7873, -2166, 7925, 1974, -7973, -1784, 8015, 1590, -8054, -1398, 8087, 1203, -8116, -1010, 8140, 814, -8160, -620, 8174, 424, -8185, -230, 
--8189, 34, -8191, 160, 8186, -356, -8179, 549, 8165, -744, -8148, 936, 8125, -1130, -8099, 1320, 8067, -1512, -8032, 1701, 7991, -1890, -7948, 2076, 7898, -2263, -7846, 2447, 7787, -2631, 
---7726, 2811, 7659, -2991, -7590, 3168, 7515, -3345, -7438, 3518, 7355, -3691, -7270, 3859, 7179, -4027, -7086, 4191, 6987, -4355, -6887, 4514, 6782, -4672, -6674, 4826, 6561, -4979, -6447, 5127, 
--6328, -5274, -6207, 5416, 6081, -5557, -5954, 5693, 5822, -5828, -5689, 5958, 5551, -6087, -5412, 6210, 5269, -6331, -5125, 6448, 4976, -6563, -4828, 6672, 4674, -6779, -4521, 6881, 4363, -6982, 
---4205, 7076, 4043, -7169, -3881, 7256, 3716, -7342, -3550, 7421, 3381, -7499, -3213, 7570, 3041, -7640, -2870, 7703, 2695, -7765, -2521, 7821, 2344, -7875, -2168, 7922, 1989, -7968, -1812, 8008, 
--1631, -8045, -1453, 8076, 1271, -8106, -1091, 8129, 909, -8150, -728, 8166, 546, -8179, -365, 8186, 182, -8191, -1, 8190, -181, -8187, 361, 8178, -543, -8167, 722, 8150, -903, -8131, 
--1081, 8106, -1261, -8080, 1437, 8047, -1615, -8013, 1790, 7972, -1965, -7930, 2138, 7883, -2311, -7833, 2481, 7778, -2652, -7721, 2819, 7659, -2987, -7595, 3151, 7525, -3316, -7454, 3476, 7378, 
---3637, -7300, 3794, 7217, -3951, -7133, 4105, 7043, -4258, -6952, 4406, 6856, -4555, -6759, 4699, 6657, -4843, -6554, 4983, 6446, -5122, -6338, 5257, 6224, -5391, -6110, 5520, 5991, -5649, -5872, 
--5773, 5748, -5897, -5623, 6015, 5494, -6133, -5365, 6246, 5232, -6358, -5098, 6465, 4960, -6570, -4823, 6671, 4681, -6771, -4539, 6866, 4393, -6959, -4248, 7047, 4099, -7134, -3950, 7216, 3798, 
---7297, -3646, 7372, 3491, -7446, -3336, 7515, 3179, -7582, -3022, 7644, 2861, -7705, -2702, 7760, 2540, -7813, -2379, 7862, 2215, -7909, -2052, 7950, 1887, -7990, -1723, 8025, 1556, -8058, -1391, 
--8085, 1224, -8112, -1058, 8132, 890, -8152, -724, 8165, 556, -8178, -390, 8185, 221, -8190, -55, 8190, -113, -8189, 278, 8182, -446, -8174, 611, 8161, -777, -8146, 942, 8126, -1107, 
---8105, 1270, 8078, -1434, -8050, 1595, 8017, -1758, -7983, 1917, 7943, -2078, -7902, 2236, 7857, -2394, -7810, 2550, 7758, -2706, -7704, 2859, 7646, -3012, -7587, 3162, 7523, -3313, -7458, 3460, 
--7389, -3608, -7318, 3752, 7243, -3897, -7167, 4038, 7086, -4179, -7004, 4316, 6918, -4453, -6831, 4587, 6740, -4720, -6648, 4850, 6552, -4979, -6456, 5105, 6355, -5230, -6253, 5351, 6148, -5472, 
---6042, 5589, 5932, -5706, -5822, 5818, 5708, -5930, -5594, 6037, 5476, -6144, -5358, 6247, 5236, -6349, -5115, 6447, 4989, -6544, -4864, 6637, 4735, -6729, -4607, 6816, 4475, -6903, -4344, 6985, 
--4209, -7067, -4075, 7144, 3938, -7220, -3801, 7291, 3661, -7362, -3522, 7428, 3380, -7493, -3239, 7554, 3094, -7613, -2951, 7668, 2805, -7722, -2660, 7771, 2513, -7820, -2367, 7863, 2218, -7906, 
---2070, 7944, 1920, -7981, -1772, 8013, 1621, -8044, -1471, 8071, 1320, -8096, -1170, 8117, 1018, -8137, -867, 8152, 715, -8166, -565, 8176, 412, -8185, -262, 8188, 110, -8191, 41, 8190, 
---192, -8187, 342, 8180, -493, -8172, 642, 8159, -793, -8145, 941, 8127, -1091, -8108, 1238, 8085, -1386, -8061, 1532, 8032, -1679, -8002, 1823, 7968, -1969, -7933, 2111, 7894, -2255, -7854, 
--2396, 7810, -2538, -7765, 2677, 7716, -2817, -7667, 2953, 7613, -3091, -7558, 3225, 7499, -3361, -7440, 3493, 7377, -3625, -7313, 3755, 7245, -3885, -7177, 4011, 7105, -4138, -7033, 4262, 6956, 
---4386, -6880, 4507, 6799, -4628, -6718, 4745, 6634, -4863, -6549, 4977, 6461, -5092, -6372, 5202, 6280, -5313, -6188, 5420, 6092, -5528, -5997, 5631, 5898, -5735, -5799, 5835, 5697, -5935, -5595, 
--6031, 5489, -6127, -5384, 6219, 5276, -6311, -5168, 6399, 5056, -6487, -4946, 6571, 4832, -6655, -4719, 6735, 4602, -6815, -4487, 6891, 4368, -6966, -4250, 7038, 4129, -7109, -4009, 7176, 3886, 
---7243, -3764, 7306, 3639, -7369, -3516, 7427, 3389, -7486, -3264, 7540, 3136, -7593, -3009, 7643, 2880, -7692, -2752, 7737, 2621, -7782, -2492, 7823, 2360, -7863, -2230, 7900, 2097, -7935, -1966, 
--7967, 1833, -7999, -1702, 8026, 1568, -8053, -1435, 8075, 1301, -8098, -1169, 8116, 1034, -8134, -901, 8148, 767, -8162, -634, 8171, 499, -8180, -366, 8185, 232, -8190, -99, 8190, -35, 
---8191, 167, 8187, -301, -8183, 432, 8175, -566, -8167, 697, 8155, -829, -8143, 959, 8126, -1091, -8110, 1220, 8089, -1351, -8068, 1479, 8044, -1608, -8019, 1735, 7990, -1864, -7962, 1989, 
--7929, -2116, -7896, 2241, 7860, -2366, -7824, 2489, 7783, -2613, -7743, 2734, 7699, -2856, -7655, 2975, 7607, -3096, -7560, 3213, 7508, -3332, -7457, 3447, 7402, -3564, -7348, 3677, 7290, -3791, 
---7232, 3903, 7170, -4015, -7109, 4124, 7044, -4234, -6980, 4340, 6912, -4448, -6845, 4552, 6774, -4657, -6703, 4759, 6629, -4861, -6556, 4961, 6479, -5060, -6403, 5157, 6323, -5254, -6245, 5348, 
--6162, -5443, -6081, 5534, 5996, -5625, -5912, 5713, 5825, -5802, -5739, 5888, 5649, -5973, -5561, 6056, 5469, -6139, -5378, 6218, 5284, -6298, -5191, 6374, 5095, -6451, -5000, 6524, 4903, -6598, 
---4806, 6668, 4706, -6739, -4608, 6806, 4506, -6873, -4406, 6937, 4303, -7001, -4202, 7062, 4097, -7123, -3994, 7180, 3888, -7238, -3784, 7292, 3677, -7346, -3571, 7397, 3463, -7448, -3356, 7496, 
--3246, -7544, -3139, 7588, 3028, -7633, -2919, 7674, 2808, -7715, -2699, 7752, 2587, -7790, -2476, 7825, 2364, -7859, -2253, 7891, 2140, -7922, -2028, 7950, 1915, -7978, -1803, 8002, 1689, -8027, 
---1577, 8048, 1463, -8070, -1350, 8088, 1236, -8106, -1123, 8121, 1009, -8136, -896, 8147, 782, -8159, -670, 8168, 555, -8176, -443, 8181, 329, -8187, -217, 8189, 103, -8191, 9, 8190, 
---122, -8190, 233, 8185, -346, -8182, 457, 8174, -570, -8168, 680, 8157, -792, -8148, 901, 8134, -1012, -8122, 1121, 8106, -1232, -8090, 1339, 8071, -1449, -8053, 1556, 8031, -1665, -8009, 
--1771, 7985, -1878, -7961, 1983, 7933, -2090, -7906, 2194, 7876, -2299, -7847, 2402, 7814, -2506, -7782, 2608, 7747, -2711, -7712, 2811, 7674, -2913, -7637, 3011, 7597, -3112, -7557, 3209, 7514, 
---3308, -7472, 3404, 7427, -3501, -7383, 3596, 7335, -3691, -7289, 3784, 7239, -3879, -7190, 3970, 7138, -4062, -7087, 4152, 7033, -4243, -6980, 4331, 6924, -4420, -6869, 4506, 6811, -4594, -6753, 
--4678, 6693, -4763, -6634, 4846, 6572, -4930, -6511, 5010, 6447, -5092, -6385, 5171, 6319, -5251, -6255, 5328, 6187, -5406, -6121, 5481, 6052, -5557, -5984, 5630, 5914, -5704, -5845, 5775, 5773, 
---5847, -5702, 5915, 5628, -5985, -5556, 6052, 5481, -6120, -5408, 6185, 5331, -6251, -5257, 6313, 5179, -6377, -5103, 6438, 5024, -6499, -4947, 6558, 4867, -6617, -4789, 6673, 4708, -6731, -4629, 
--6785, 4547, -6840, -4467, 6892, 4384, -6945, -4303, 6995, 4219, -7046, -4137, 7094, 4052, -7142, -3970, 7188, 3884, -7234, -3801, 7278, 3715, -7322, -3630, 7363, 3544, -7405, -3459, 7445, 3372, 
---7485, -3286, 7521, 3198, -7559, -3112, 7594, 3024, -7630, -2938, 7662, 2849, -7696, -2762, 7726, 2673, -7758, -2586, 7786, 2497, -7816, -2409, 7842, 2320, -7869, -2232, 7893, 2143, -7918, -2055, 
--7940, 1965, -7963, -1877, 7983, 1787, -8004, -1699, 8022, 1609, -8041, -1521, 8056, 1431, -8073, -1343, 8087, 1253, -8102, -1165, 8114, 1075, -8126, -987, 8136, 897, -8147, -810, 8155, 720, 
---8164, -633, 8169, 543, -8176, -456, 8180, 367, -8185, -280, 8187, 192, -8190, -105, 8190, 17, -8191, 69, 8190, -157, -8189, 243, 8185, -331, -8183, 416, 8178, -503, -8173, 588, 
--8166, -674, -8160, 758, 8151, -844, -8143, 928, 8133, -1014, -8123, 1097, 8111, -1181, -8100, 1264, 8086, -1348, -8073, 1430, 8057, -1513, -8043, 1594, 8026, -1677, -8009, 1757, 7991, -1839, 
---7973, 1919, 7953, -2000, -7933, 2079, 7912, -2159, -7891, 2238, 7868, -2317, -7845, 2394, 7821, -2473, -7797, 2549, 7771, -2627, -7746, 2703, 7718, -2780, -7692, 2854, 7663, -2930, -7635, 3004, 
--7605, -3079, -7576, 3152, 7544, -3226, -7514, 3298, 7481, -3371, -7450, 3442, 7415, -3514, -7383, 3584, 7347, -3655, -7314, 3724, 7277, -3794, -7242, 3862, 7204, -3931, -7168, 3997, 7130, -4066, 
---7092, 4131, 7053, -4198, -7014, 4263, 6974, -4329, -6934, 4392, 6893, -4457, -6852, 4519, 6810, -4583, -6768, 4644, 6725, -4707, -6683, 4767, 6638, -4829, -6595, 4888, 6550, -4948, -6506, 5006, 
--6460, -5066, -6415, 5122, 6368, -5180, -6322, 5236, 6274, -5293, -6228, 5348, 6180, -5404, -6133, 5457, 6083, -5512, -6036, 5564, 5986, -5617, -5938, 5668, 5887, -5721, -5838, 5771, 5787, -5822, 
---5737, 5871, 5685, -5921, -5635, 5969, 5583, -6018, -5532, 6064, 5479, -6112, -5428, 6157, 5375, -6204, -5323, 6248, 5269, -6293, -5217, 6336, 5163, -6381, -5110, 6423, 5056, -6466, -5003, 6507, 
--4947, -6549, -4894, 6588, 4839, -6629, -4785, 6668, 4729, -6707, -4675, 6745, 4619, -6783, -4565, 6819, 4508, -6857, -4454, 6892, 4397, -6929, -4342, 6962, 4285, -6998, -4230, 7031, 4173, -7065, 
---4118, 7097, 4061, -7130, -4005, 7160, 3948, -7193, -3892, 7222, 3835, -7253, -3779, 7282, 3721, -7312, -3666, 7339, 3608, -7368, -3552, 7394, 3494, -7422, -3438, 7447, 3380, -7474, -3324, 7498, 
--3266, -7524, -3210, 7548, 3152, -7572, -3096, 7595, 3038, -7618, -2982, 7640, 2924, -7662, -2868, 7683, 2811, -7704, -2755, 7724, 2697, -7744, -2641, 7763, 2583, -7783, -2528, 7800, 2470, -7819, 
---2414, 7835, 2357, -7853, -2301, 7869, 2244, -7886, -2189, 7901, 2132, -7917, -2076, 7930, 2019, -7946, -1964, 7958, 1908, -7973, -1853, 7985, 1796, -7998, -1742, 8009, 1685, -8022, -1631, 8032, 
--1575, -8044, -1520, 8053, 1464, -8064, -1411, 8073, 1355, -8083, -1301, 8091, 1246, -8100, -1192, 8107, 1137, -8116, -1084, 8122, 1029, -8130, -977, 8135, 922, -8142, -870, 8147, 815, -8153, 
---763, 8157, 709, -8163, -657, 8166, 604, -8171, -552, 8174, 499, -8178, -448, 8180, 395, -8183, -344, 8184, 292, -8187, -242, 8188, 189, -8190, -139, 8190, 88, -8191, -38, 8190, 
---13, -8191, 63, 8190, -114, -8190, 162, 8188, -213, -8188, 261, 8185, -312, -8185, 360, 8181, -409, -8180, 457, 8176, -506, -8174, 553, 8170, -602, -8168, 649, 8163, -698, -8160, 
--744, 8154, -792, -8151, 838, 8145, -885, -8141, 931, 8135, -978, -8130, 1023, 8123, -1069, -8118, 1114, 8111, -1160, -8106, 1204, 8098, -1250, -8092, 1293, 8084, -1339, -8078, 1382, 8069, 
---1427, -8063, 1469, 8054, -1514, -8046, 1556, 8037, -1600, -8030, 1641, 8020, -1685, -8012, 1726, 8002, -1769, -7994, 1809, 7983, -1852, -7975, 1892, 7964, -1934, -7955, 1974, 7944, -2015, -7935, 
--2054, 7923, -2095, -7914, 2134, 7902, -2175, -7892, 2213, 7880, -2253, -7870, 2291, 7858, -2330, -7847, 2368, 7835, -2407, -7824, 2443, 7812, -2482, -7801, 2518, 7788, -2556, -7776, 2592, 7763, 
---2630, -7752, 2665, 7738, -2702, -7727, 2737, 7713, -2773, -7701, 2808, 7688, -2844, -7676, 2878, 7662, -2913, -7649, 2947, 7635, -2982, -7623, 3015, 7609, -3049, -7596, 3082, 7582, -3116, -7569, 
--3148, 7554, -3182, -7542, 3213, 7527, -3246, -7514, 3277, 7499, -3310, -7486, 3340, 7471, -3373, -7458, 3403, 7443, -3434, -7430, 3464, 7415, -3495, -7401, 3524, 7386, -3555, -7373, 3584, 7358, 
---3614, -7344, 3642, 7329, -3672, -7315, 3700, 7300, -3729, -7286, 3756, 7271, -3785, -7257, 3812, 7242, -3840, -7228, 3867, 7213, -3895, -7199, 3920, 7184, -3948, -7170, 3973, 7155, -4000, -7141, 
--4025, 7126, -4052, -7112, 4076, 7096, -4103, -7083, 4127, 7067, -4153, -7054, 4176, 7038, -4201, -7025, 4225, 7009, -4249, -6996, 4272, 6981, -4297, -6967, 4319, 6952, -4343, -6939, 4365, 6923, 
---4388, -6910, 4410, 6895, -4433, -6881, 4454, 6866, -4477, -6853, 4497, 6838, -4520, -6825, 4540, 6810, -4562, -6797, 4581, 6782, -4603, -6769, 4622, 6754, -4643, -6742, 4662, 6727, -4683, -6714, 
--4701, 6700, -4722, -6687, 4740, 6673, -4760, -6660, 4778, 6646, -4797, -6634, 4814, 6619, -4833, -6607, 4850, 6593, -4869, -6581, 4886, 6567, -4904, -6555, 4920, 6541, -4938, -6530, 4954, 6516, 
---4971, -6504, 4987, 6491, -5004, -6479, 5019, 6466, -5036, -6455, 5051, 6442, -5067, -6431, 5081, 6418, -5097, -6407, 5111, 6394, -5127, -6383, 5141, 6370, -5156, -6360, 5169, 6347, -5184, -6337, 
--5197, 6325, -5212, -6314, 5224, 6302, -5238, -6292, 5251, 6280, -5265, -6271, 5276, 6259, -5290, -6249, 5301, 6238, -5315, -6228, 5326, 6217, -5339, -6208, 5349, 6197, -5362, -6188, 5372, 6177, 
---5385, -6168, 5395, 6158, -5407, -6149, 5417, 6139, -5428, -6130, 5438, 6120, -5449, -6112, 5458, 6102, -5469, -6094, 5478, 6085, -5488, -6077, 5497, 6068, -5507, -6060, 5515, 6051, -5525, -6044, 
--5533, 6035, -5543, -6028, 5550, 6019, -5560, -6012, 5567, 6004, -5576, -5997, 5583, 5989, -5591, -5983, 5598, 5975, -5607, -5969, 5613, 5961, -5621, -5956, 5627, 5948, -5635, -5943, 5640, 5935, 
---5648, -5930, 5653, 5923, -5661, -5918, 5666, 5912, -5673, -5907, 5677, 5900, -5684, -5896, 5689, 5890, -5695, -5886, 5699, 5880, -5705, -5876, 5709, 5870, -5715, -5867, 5718, 5861, -5724, -5858, 
--5727, 5853, -5732, -5850, 5736, 5845, -5740, -5842, 5743, 5837, -5748, -5835, 5750, 5831, -5755, -5828, 5757, 5824, -5761, -5822, 5763, 5819, -5767, -5817, 5768, 5813, -5772, -5812, 5773, 5809, 
---5776, -5808, 5777, 5805, -5780, -5804, 5781, 5801, -5784, -5800, 5784, 5798, -5786, -5798, 5787, 5796, -5789, -5796, 5789, 5794, -5790, -5794, 5790, 5792, -5792, -5793, 5791, 5792, -5792, -5792, 
--5791, 5791, -5792, -5793, 5791, 5792, -5792, -5793, 5790, 5793, -5791, -5794, 5789, 5794, -5789, -5796, 5787, 5796, -5787, -5798, 5785, 5799, -5784, -5801, 5782, 5802, -5781, -5805, 5778, 5806, 
---5777, -5809, 5774, 5810, -5773, -5813, 5769, 5815, -5768, -5818, 5764, 5820, -5762, -5824, 5758, 5826, -5756, -5830, 5752, 5832, -5750, -5837, 5745, 5839, -5742, -5844, 5738, 5847, -5735, -5852, 
--5729, 5855, -5726, -5860, 5721, 5863, -5717, -5869, 5712, 5873, -5708, -5878, 5702, 5882, -5698, -5888, 5691, 5892, -5687, -5899, 5680, 5903, -5676, -5910, 5669, 5914, -5664, -5921, 5657, 5926, 
---5651, -5933, 5644, 5939, -5638, -5946, 5630, 5951, -5624, -5959, 5616, 5965, -5610, -5973, 5602, 5978, -5595, -5987, 5587, 5993, -5580, -6001, 5571, 6008, -5564, -6016, 5554, 6023, -5547, -6032, 
--5537, 6039, -5530, -6048, 5520, 6055, -5512, -6064, 5501, 6072, -5493, -6081, 5482, 6089, -5474, -6099, 5463, 6107, -5454, -6117, 5443, 6125, -5433, -6135, 5422, 6143, -5412, -6154, 5400, 6163, 
---5390, -6173, 5378, 6182, -5368, -6193, 5355, 6202, -5345, -6213, 5332, 6222, -5321, -6234, 5308, 6243, -5296, -6255, 5283, 6264, -5271, -6276, 5257, 6286, -5245, -6298, 5231, 6308, -5218, -6320, 
--5204, 6330, -5191, -6343, 5176, 6353, -5163, -6366, 5148, 6376, -5134, -6389, 5119, 6400, -5105, -6413, 5089, 6424, -5075, -6437, 5058, 6448, -5044, -6461, 5027, 6472, -5012, -6486, 4995, 6497, 
---4980, -6511, 4962, 6522, -4947, -6536, 4929, 6548, -4913, -6562, 4894, 6574, -4878, -6588, 4859, 6600, -4842, -6614, 4823, 6626, -4806, -6640, 4787, 6653, -4769, -6667, 4749, 6679, -4731, -6694, 
--4711, 6706, -4693, -6721, 4672, 6734, -4653, -6749, 4632, 6761, -4613, -6776, 4592, 6789, -4572, -6804, 4550, 6817, -4530, -6832, 4508, 6845, -4488, -6860, 4465, 6873, -4444, -6889, 4421, 6902, 
---4400, -6917, 4376, 6930, -4354, -6946, 4330, 6959, -4308, -6974, 4284, 6988, -4261, -7003, 4237, 7017, -4214, -7032, 4188, 7046, -4165, -7061, 4139, 7075, -4115, -7090, 4089, 7104, -4065, -7119, 
--4038, 7133, -4013, -7148, 3986, 7162, -3961, -7178, 3934, 7191, -3908, -7207, 3880, 7220, -3854, -7236, 3826, 7249, -3799, -7265, 3770, 7278, -3743, -7294, 3714, 7307, -3686, -7323, 3657, 7336, 
---3629, -7351, 3598, 7365, -3570, -7380, 3539, 7393, -3510, -7409, 3479, 7422, -3450, -7437, 3418, 7450, -3388, -7465, 3356, 7478, -3326, -7493, 3293, 7506, -3262, -7521, 3229, 7534, -3198, -7549, 
--3164, 7561, -3132, -7576, 3098, 7588, -3066, -7603, 3032, 7615, -2999, -7630, 2964, 7642, -2931, -7656, 2895, 7668, -2861, -7682, 2825, 7694, -2791, -7708, 2755, 7720, -2720, -7733, 2683, 7745, 
---2648, -7758, 2610, 7769, -2575, -7783, 2537, 7794, -2501, -7807, 2462, 7817, -2426, -7830, 2387, 7841, -2349, -7853, 2310, 7864, -2272, -7876, 2232, 7886, -2194, -7898, 2154, 7907, -2115, -7919, 
--2074, 7929, -2035, -7940, 1994, 7949, -1954, -7960, 1913, 7969, -1873, -7980, 1830, 7988, -1790, -7998, 1747, 8007, -1706, -8016, 1662, 8024, -1621, -8034, 1577, 8041, -1535, -8051, 1491, 8058, 
---1448, -8066, 1404, 8073, -1361, -8081, 1316, 8088, -1272, -8096, 1227, 8101, -1183, -8109, 1137, 8114, -1092, -8121, 1046, 8126, -1001, -8133, 954, 8137, -909, -8144, 861, 8148, -815, -8153, 
--767, 8157, -721, -8162, 673, 8165, -626, -8169, 577, 8172, -530, -8176, 481, 8178, -434, -8181, 384, 8183, -336, -8186, 286, 8186, -238, -8189, 187, 8189, -139, -8191, 88, 8190, 
---39, -8191, -13, 8190, 62, -8191, -114, 8189, 164, -8189, -216, 8187, 266, -8186, -319, 8183, 369, -8182, -422, 8178, 473, -8176, -526, 8172, 578, -8169, -631, 8164, 683, -8161, 
---737, 8155, 789, -8151, -843, 8144, 895, -8139, -950, 8132, 1002, -8127, -1057, 8118, 1110, -8112, -1165, 8103, 1219, -8096, -1274, 8087, 1328, -8079, -1383, 8068, 1437, -8059, -1493, 8048, 
--1547, -8039, -1603, 8027, 1657, -8016, -1714, 8003, 1768, -7992, -1825, 7978, 1880, -7966, -1936, 7952, 1991, -7939, -2048, 7923, 2104, -7909, -2161, 7893, 2216, -7878, -2273, 7861, 2329, -7845, 
---2386, 7827, 2442, -7810, -2499, 7791, 2555, -7773, -2613, 7753, 2668, -7735, -2726, 7714, 2782, -7694, -2840, 7672, 2896, -7651, -2954, 7628, 3010, -7607, -3068, 7583, 3124, -7560, -3182, 7535, 
--3238, -7512, -3296, 7486, 3352, -7461, -3410, 7434, 3466, -7409, -3523, 7381, 3579, -7354, -3637, 7325, 3693, -7297, -3751, 7267, 3806, -7238, -3864, 7207, 3920, -7177, -3977, 7145, 4033, -7114, 
---4090, 7080, 4145, -7048, -4202, 7014, 4257, -6981, -4314, 6945, 4369, -6911, -4426, 6874, 4481, -6839, -4537, 6801, 4591, -6765, -4648, 6726, 4702, -6688, -4758, 6648, 4811, -6609, -4867, 6568, 
--4920, -6528, -4976, 6486, 5029, -6445, -5083, 6401, 5136, -6359, -5191, 6314, 5243, -6271, -5297, 6225, 5349, -6181, -5402, 6134, 5453, -6088, -5506, 6040, 5557, -5994, -5610, 5944, 5660, -5896, 
---5712, 5846, 5762, -5797, -5813, 5745, 5862, -5695, -5913, 5643, 5961, -5591, -6011, 5537, 6059, -5485, -6109, 5430, 6156, -5376, -6205, 5320, 6251, -5265, -6299, 5208, 6345, -5152, -6392, 5093, 
--6437, -5036, -6483, 4977, 6527, -4919, -6573, 4858, 6616, -4799, -6661, 4737, 6703, -4676, -6747, 4613, 6789, -4552, -6832, 4488, 6872, -4425, -6914, 4360, 6954, -4296, -6995, 4230, 7033, -4165, 
---7073, 4098, 7111, -4032, -7150, 3964, 7186, -3897, -7224, 3827, 7259, -3759, -7296, 3689, 7330, -3620, -7366, 3548, 7399, -3478, -7433, 3406, 7465, -3335, -7498, 3262, 7529, -3190, -7561, 3115, 
--7590, -3042, -7621, 2967, 7649, -2893, -7678, 2817, 7705, -2742, -7733, 2665, 7758, -2589, -7784, 2511, 7808, -2434, -7834, 2355, 7856, -2278, -7880, 2198, 7901, -2120, -7923, 2039, 7943, -1960, 
---7963, 1879, 7981, -1799, -8001, 1717, 8017, -1636, -8035, 1553, 8050, -1472, -8066, 1388, 8079, -1306, -8093, 1222, 8105, -1140, -8118, 1055, 8128, -971, -8139, 886, 8147, -802, -8156, 716, 
--8163, -631, -8170, 545, 8175, -460, -8181, 373, 8184, -287, -8188, 200, 8189, -114, -8191, 26, 8190, 60, -8191, -149, 8188, 236, -8187, -324, 8182, 411, -8179, -500, 8172, 588, 
---8167, -677, 8159, 765, -8151, -854, 8141, 942, -8132, -1032, 8120, 1119, -8108, -1209, 8094, 1297, -8081, -1387, 8064, 1475, -8049, -1565, 8031, 1653, -8013, -1743, 7993, 1831, -7974, -1921, 
--7951, 2009, -7930, -2099, 7905, 2187, -7882, -2277, 7855, 2364, -7829, -2454, 7800, 2541, -7773, -2630, 7742, 2717, -7712, -2806, 7679, 2893, -7647, -2981, 7612, 3068, -7577, -3156, 7540, 3242, 
---7504, -3329, 7464, 3415, -7426, -3502, 7384, 3587, -7343, -3673, 7300, 3757, -7257, -3843, 7211, 3926, -7166, -4012, 7118, 4094, -7070, -4179, 7020, 4260, -6971, -4344, 6918, 4425, -6867, -4507, 
--6812, 4588, -6758, -4669, 6702, 4748, -6646, -4829, 6587, 4907, -6529, -4986, 6468, 5063, -6408, -5142, 6345, 5217, -6283, -5295, 6217, 5369, -6153, -5445, 6086, 5518, -6019, -5593, 5950, 5665, 
---5882, -5738, 5810, 5808, -5740, -5880, 5666, 5949, -5594, -6019, 5518, 6086, -5444, -6155, 5366, 6221, -5290, -6287, 5211, 6351, -5132, -6417, 5051, 6479, -4971, -6542, 4888, 6603, -4805, -6664, 
--4720, 6723, -4636, -6783, 4549, 6839, -4464, -6897, 4375, 6952, -4288, -7007, 4197, 7060, -4108, -7113, 4016, 7164, -3925, -7215, 3831, 7264, -3739, -7313, 3643, 7359, -3549, -7406, 3452, 7449, 
---3357, -7494, 3258, 7535, -3161, -7578, 3061, 7617, -2963, -7656, 2861, 7693, -2761, -7730, 2659, 7764, -2558, -7799, 2454, 7830, -2351, -7862, 2246, 7891, -2142, -7921, 2036, 7947, -1931, -7973, 
--1824, 7997, -1718, -8021, 1610, 8041, -1503, -8062, 1394, 8080, -1286, -8098, 1176, 8113, -1067, -8129, 956, 8141, -847, -8153, 735, 8162, -625, -8172, 513, 8178, -402, -8184, 289, 8187, 
---178, -8191, 65, 8190, 47, -8191, -160, 8188, 272, -8185, -386, 8179, 499, -8173, -613, 8163, 725, -8154, -840, 8141, 952, -8129, -1067, 8113, 1179, -8098, -1294, 8079, 1406, -8060, 
---1520, 8037, 1632, -8015, -1747, 7990, 1858, -7964, -1972, 7935, 2084, -7907, -2197, 7875, 2308, -7843, -2421, 7807, 2531, -7772, -2643, 7733, 2753, -7695, -2864, 7653, 2973, -7611, -3084, 7566, 
--3192, -7520, -3302, 7472, 3409, -7423, -3517, 7371, 3623, -7320, -3731, 7264, 3836, -7210, -3942, 7151, 4045, -7093, -4150, 7031, 4252, -6970, -4355, 6905, 4456, -6840, -4558, 6772, 4657, -6704, 
---4757, 6633, 4854, -6562, -4952, 6487, 5048, -6413, -5144, 6336, 5237, -6259, -5332, 6178, 5423, -6098, -5515, 6014, 5605, -5931, -5695, 5845, 5782, -5759, -5869, 5669, 5954, -5580, -6039, 5488, 
--6121, -5396, -6204, 5301, 6284, -5206, -6364, 5108, 6441, -5011, -6518, 4911, 6592, -4811, -6667, 4708, 6738, -4605, -6810, 4500, 6878, -4395, -6947, 4287, 7012, -4179, -7077, 4069, 7139, -3959, 
---7202, 3847, 7260, -3735, -7320, 3620, 7375, -3506, -7431, 3389, 7483, -3273, -7535, 3154, 7583, -3036, -7632, 2915, 7677, -2795, -7722, 2673, 7763, -2551, -7804, 2427, 7841, -2304, -7879, 2178, 
--7913, -2053, -7946, 1926, 7976, -1800, -8005, 1671, 8031, -1544, -8057, 1414, 8078, -1286, -8100, 1155, 8118, -1026, -8135, 894, 8148, -763, -8162, 631, 8171, -500, -8180, 366, 8185, -234, 
---8190, 101, 8190, 32, -8191, -166, 8187, 299, -8183, -433, 8175, 566, -8167, -701, 8155, 833, -8142, -968, 8125, 1101, -8108, -1235, 8086, 1368, -8065, -1502, 8039, 1634, -8013, -1768, 
--7983, 1899, -7952, -2033, 7917, 2163, -7882, -2296, 7843, 2426, -7803, -2557, 7760, 2686, -7716, -2816, 7667, 2944, -7619, -3073, 7566, 3199, -7513, -3327, 7456, 3452, -7399, -3578, 7337, 3701, 
---7276, -3826, 7210, 3947, -7144, -4070, 7073, 4189, -7003, -4310, 6928, 4427, -6854, -4545, 6775, 4660, -6696, -4776, 6613, 4889, -6530, -5002, 6443, 5112, -6356, -5222, 6265, 5330, -6174, -5437, 
--6079, 5542, -5984, -5646, 5885, 5748, -5786, -5849, 5683, 5947, -5580, -6045, 5474, 6140, -5368, -6235, 5257, 6326, -5148, -6417, 5034, 6505, -4921, -6592, 4804, 6676, -4687, -6759, 4567, 6839, 
---4447, -6919, 4324, 6994, -4201, -7070, 4074, 7141, -3949, -7212, 3819, 7279, -3691, -7346, 3559, 7408, -3427, -7471, 3293, 7529, -3159, -7586, 3022, 7639, -2886, -7692, 2746, 7741, -2608, -7789, 
--2467, 7832, -2326, -7875, 2183, 7914, -2041, -7952, 1896, 7985, -1752, -8018, 1605, 8046, -1460, -8073, 1311, 8096, -1165, -8119, 1015, 8136, -868, -8153, 717, 8165, -568, -8177, 417, 8183, 
---268, -8189, 116, 8190, 34, -8191, -186, 8186, 336, -8181, -489, 8171, 639, -8160, -792, 8144, 942, -8128, -1094, 8107, 1244, -8084, -1396, 8057, 1546, -8029, -1697, 7997, 1846, -7963, 
---1996, 7925, 2144, -7885, -2293, 7841, 2439, -7796, -2587, 7747, 2732, -7696, -2879, 7641, 3022, -7584, -3167, 7523, 3309, -7461, -3451, 7395, 3591, -7328, -3732, 7256, 3869, -7183, -4007, 7105, 
--4142, -7027, -4277, 6944, 4409, -6861, -4542, 6772, 4671, -6684, -4800, 6590, 4926, -6496, -5053, 6398, 5175, -6299, -5298, 6195, 5417, -6092, -5536, 5983, 5651, -5875, -5766, 5762, 5877, -5648, 
---5988, 5530, 6095, -5413, -6201, 5290, 6304, -5168, -6406, 5042, 6504, -4915, -6601, 4785, 6694, -4654, -6787, 4520, 6875, -4385, -6962, 4247, 7045, -4109, -7127, 3967, 7204, -3825, -7281, 3680, 
--7353, -3535, -7424, 3387, 7491, -3238, -7556, 3087, 7617, -2936, -7676, 2782, 7731, -2628, -7784, 2472, 7833, -2316, -7880, 2157, 7923, -1998, -7964, 1837, 8000, -1677, -8035, 1514, 8064, -1353, 
---8092, 1188, 8115, -1025, -8137, 859, 8154, -695, -8169, 528, 8178, -363, -8187, 195, 8190, -29, -8191, -139, 8187, 305, -8182, -473, 8172, 640, -8159, -808, 8142, 974, -8123, -1142, 
--8098, 1307, -8073, -1474, 8041, 1639, -8008, -1806, 7970, 1969, -7930, -2134, 7885, 2297, -7839, -2460, 7787, 2621, -7733, -2782, 7674, 2941, -7614, -3101, 7548, 3257, -7481, -3414, 7409, 3568, 
---7335, -3723, 7257, 3874, -7176, -4025, 7091, 4173, -7004, -4321, 6912, 4466, -6819, -4611, 6721, 4751, -6622, -4892, 6517, 5029, -6412, -5166, 6302, 5298, -6190, -5431, 6074, 5559, -5957, -5686, 
--5835, 5809, -5712, -5932, 5585, 6050, -5456, -6168, 5324, 6281, -5190, -6393, 5052, 6500, -4914, -6607, 4771, 6708, -4628, -6809, 4480, 6904, -4333, -6998, 4181, 7088, -4029, -7176, 3873, 7258, 
---3717, -7340, 3557, 7416, -3397, -7491, 3233, 7560, -3070, -7628, 2903, 7690, -2736, -7750, 2567, 7805, -2397, -7859, 2224, 7906, -2052, -7952, 1877, 7992, -1703, -8031, 1526, 8063, -1350, -8094, 
--1171, 8119, -993, -8142, 812, 8159, -633, -8174, 452, 8183, -272, -8190, 89, 8190, 91, -8189, -274, 8182, 455, -8173, -637, 8158, 818, -8141, -1001, 8118, 1181, -8092, -1362, 8061, 
--1542, -8027, -1722, 7988, 1900, -7946, -2079, 7898, 2256, -7849, -2433, 7793, 2608, -7735, -2783, 7672, 2955, -7606, -3128, 7534, 3297, -7461, -3467, 7381, 3633, -7300, -3799, 7213, 3962, -7124, 
---4125, 7029, 4284, -6933, -4442, 6830, 4597, -6727, -4752, 6617, 4902, -6506, -5052, 6390, 5197, -6272, -5341, 6148, 5481, -6023, -5621, 5893, 5755, -5762, -5889, 5625, 6017, -5488, -6145, 5345, 
--6267, -5201, -6388, 5052, 6504, -4903, -6619, 4749, 6728, -4594, -6835, 4434, 6937, -4274, -7038, 4109, 7132, -3944, -7225, 3775, 7312, -3605, -7397, 3431, 7477, -3257, -7554, 3080, 7625, -2902, 
---7694, 2720, 7757, -2539, -7817, 2355, 7872, -2170, -7924, 1983, 7970, -1796, -8013, 1606, 8050, -1417, -8084, 1225, 8112, -1034, -8138, 840, 8157, -647, -8173, 452, 8183, -259, -8190, 63, 
--8190, 131, -8188, -327, 8180, 521, -8168, -718, 8150, 911, -8129, -1107, 8102, 1300, -8071, -1495, 8035, 1687, -7995, -1880, 7949, 2070, -7900, -2261, 7845, 2449, -7787, -2638, 7722, 2823, 
---7655, -3010, 7581, 3192, -7505, -3375, 7422, 3554, -7337, -3733, 7245, 3908, -7151, -4083, 7051, 4253, -6948, -4424, 6839, 4589, -6728, -4755, 6611, 4915, -6492, -5075, 6367, 5230, -6239, -5384, 
--6106, 5533, -5972, -5680, 5831, 5823, -5689, -5964, 5541, 6099, -5392, -6233, 5237, 6361, -5081, -6488, 4920, 6609, -4757, -6727, 4589, 6840, -4421, -6951, 4247, 7055, -4073, -7157, 3894, 7253, 
---3715, -7347, 3531, 7434, -3346, -7518, 3158, 7596, -2969, -7671, 2776, 7740, -2584, -7805, 2387, 7864, -2191, -7920, 1991, 7969, -1792, -8015, 1589, 8054, -1387, -8090, 1183, 8119, -979, -8145, 
--772, 8163, -567, -8178, 359, 8186, -153, -8191, -56, 8189, 263, -8183, -471, 8170, 678, -8154, -886, 8131, 1092, -8104, -1300, 8070, 1505, -8032, -1711, 7987, 1914, -7939, -2118, 7884, 
--2319, -7826, -2521, 7760, 2719, -7691, -2917, 7616, 3112, -7536, -3307, 7450, 3498, -7361, -3688, 7265, 3875, -7166, -4061, 7060, 4242, -6952, -4423, 6836, 4599, -6718, -4774, 6593, 4944, -6466, 
---5113, 6332, 5277, -6196, -5439, 6053, 5596, -5908, -5751, 5757, 5900, -5604, -6047, 5445, 6188, -5285, -6328, 5118, 6461, -4950, -6591, 4776, 6716, -4601, -6838, 4420, 6953, -4238, -7065, 4051, 
--7171, -3864, -7274, 3671, 7369, -3477, -7462, 3279, 7548, -3081, -7630, 2878, 7706, -2675, -7777, 2468, 7842, -2260, -7903, 2050, 7956, -1839, -8006, 1625, 8048, -1412, -8087, 1195, 8118, -980, 
---8145, 761, 8164, -544, -8180, 324, 8188, -106, -8191, -115, 8187, 333, -8179, -554, 8164, 772, -8144, -992, 8116, 1210, -8085, -1428, 8045, 1644, -8002, -1861, 7950, 2075, -7895, -2289, 
--7832, 2500, -7766, -2712, 7691, 2919, -7613, -3127, 7527, 3330, -7438, -3533, 7341, 3732, -7240, -3930, 7132, 4124, -7021, -4316, 6902, 4504, -6780, -4690, 6651, 4871, -6518, -5050, 6379, 5224, 
---6237, -5396, 6088, 5562, -5936, -5726, 5778, 5884, -5617, -6040, 5450, 6189, -5280, -6335, 5104, 6475, -4927, -6612, 4743, 6742, -4557, -6869, 4366, 6989, -4174, -7106, 3976, 7215, -3776, -7321, 
--3572, 7419, -3367, -7514, 3157, 7601, -2946, -7684, 2731, 7759, -2516, -7830, 2296, 7893, -2077, -7952, 1853, 8003, -1630, -8050, 1404, 8088, -1178, -8122, 949, 8148, -721, -8169, 491, 8182, 
---261, -8190, 30, 8190, 200, -8185, -432, 8172, 661, -8155, -893, 8128, 1122, -8098, -1352, 8058, 1579, -8015, -1807, 7962, 2032, -7906, -2258, 7840, 2480, -7771, -2702, 7693, 2920, -7611, 
---3137, 7521, 3351, -7426, -3564, 7323, 3772, -7216, -3979, 7102, 4182, -6983, -4383, 6856, 4578, -6726, -4772, 6588, 4960, -6447, -5146, 6298, 5327, -6145, -5504, 5986, 5676, -5823, -5845, 5654, 
--6007, -5481, -6166, 5302, 6318, -5121, -6467, 4932, 6609, -4742, -6748, 4545, 6878, -4347, -7006, 4142, 7125, -3936, -7240, 3725, 7348, -3512, -7451, 3294, 7546, -3075, -7637, 2851, 7719, -2627, 
---7797, 2398, 7866, -2169, -7930, 1936, 7986, -1703, -8037, 1466, 8079, -1230, -8116, 990, 8144, -752, -8167, 511, 8181, -271, -8190, 29, 8190, 212, -8185, -455, 8170, 695, -8151, -937, 
--8122, 1176, -8088, -1417, 8045, 1654, -7997, -1892, 7940, 2127, -7878, -2362, 7807, 2593, -7731, -2824, 7645, 3051, -7556, -3277, 7457, 3499, -7353, -3719, 7241, 3934, -7125, -4148, 7000, 4357, 
---6870, -4564, 6733, 4764, -6591, -4963, 6441, 5156, -6287, -5345, 6125, 5529, -5960, -5709, 5787, 5882, -5611, -6052, 5427, 6215, -5241, -6374, 5047, 6526, -4851, -6673, 4648, 6813, -4443, -6949, 
--4231, 7076, -4018, -7199, 3798, 7313, -3577, -7423, 3351, 7524, -3123, -7620, 2890, 7707, -2656, -7789, 2418, 7861, -2179, -7929, 1936, 7987, -1692, -8040, 1446, 8083, -1199, -8121, 949, 8149, 
---701, -8171, 449, 8184, -198, -8191, -54, 8189, 305, -8180, -558, 8162, 808, -8138, -1060, 8104, 1309, -8065, -1559, 8016, 1806, -7961, -2053, 7896, 2296, -7826, -2540, 7747, 2779, -7662, 
---3018, 7567, 3251, -7467, -3484, 7358, 3712, -7243, -3939, 7120, 4159, -6991, -4378, 6853, 4591, -6711, -4801, 6560, 5005, -6405, -5206, 6241, 5401, -6073, -5592, 5897, 5776, -5717, -5956, 5529, 
--6128, -5338, -6297, 5139, 6458, -4937, -6614, 4728, 6762, -4516, -6905, 4297, 7039, -4076, -7169, 3849, 7289, -3620, -7405, 3385, 7511, -3148, -7611, 2906, 7702, -2663, -7788, 2415, 7863, -2167, 
---7933, 1914, 7993, -1661, -8047, 1404, 8091, -1147, -8128, 888, 8155, -629, -8176, 367, 8187, -106, -8191, -156, 8185, 417, -8173, -679, 8150, 939, -8121, -1201, 8082, 1459, -8036, -1718, 
--7980, 1973, -7918, -2228, 7845, 2480, -7766, -2731, 7677, 2977, -7582, -3222, 7477, 3462, -7367, -3701, 7246, 3934, -7120, -4166, 6984, 4391, -6843, -4613, 6693, 4829, -6537, -5042, 6373, 5248, 
---6203, -5450, 6025, 5645, -5843, -5836, 5652, 6019, -5457, -6198, 5254, 6368, -5047, -6534, 4833, 6690, -4616, -6842, 4391, 6985, -4164, -7122, 3929, 7250, -3693, -7372, 3450, 7484, -3206, -7590, 
--2956, 7686, -2704, -7776, 2448, 7855, -2190, -7928, 1928, 7991, -1666, -8047, 1400, 8092, -1134, -8130, 864, 8158, -596, -8179, 324, 8188, -54, -8191, -218, 8183, 488, -8168, -760, 8142, 
--1029, -8108, -1299, 8064, 1566, -8013, -1834, 7951, 2097, -7882, -2361, 7803, 2620, -7716, -2878, 7619, 3132, -7516, -3384, 7402, 3630, -7281, -3874, 7151, 4113, -7014, -4349, 6867, 4578, -6715, 
---4804, 6552, 5023, -6385, -5239, 6208, 5446, -6026, -5650, 5834, 5846, -5639, -6036, 5434, 6219, -5225, -6396, 5009, 6564, -4788, -6727, 4559, 6880, -4328, -7027, 4089, 7165, -3847, -7296, 3599, 
--7417, -3348, -7532, 3092, 7636, -2833, -7733, 2570, 7819, -2305, -7899, 2035, 7967, -1764, -8028, 1490, 8078, -1215, -8120, 937, 8152, -659, -8175, 379, 8187, -100, -8191, -181, 8184, 461, 
---8169, -742, 8143, 1020, -8109, -1300, 8063, 1576, -8010, -1852, 7946, 2124, -7873, -2396, 7790, 2664, -7699, -2930, 7597, 3191, -7488, -3451, 7368, 3704, -7241, -3955, 7103, 4200, -6959, -4442, 
--6804, 4677, -6643, -4908, 6472, 5131, -6295, -5351, 6108, 5562, -5915, -5769, 5714, 5966, -5507, -6159, 5292, 6342, -5072, -6520, 4843, 6688, -4611, -6850, 4371, 7002, -4127, -7147, 3876, 7282, 
---3623, -7409, 3362, 7526, -3099, -7636, 2831, 7734, -2560, -7825, 2285, 7904, -2008, -7976, 1727, 8035, -1445, -8087, 1159, 8127, -874, -8159, 585, 8179, -298, -8190, 8, 8189, 281, -8180, 
---571, 8159, 859, -8130, -1147, 8088, 1433, -8038, -1719, 7977, 2001, -7907, -2282, 7825, 2559, -7735, -2835, 7633, 3106, -7523, -3374, 7402, 3637, -7274, -3897, 7134, 4151, -6987, -4401, 6828, 
--4644, -6664, -4883, 6488, 5114, -6306, -5341, 6114, 5558, -5916, -5771, 5708, 5975, -5495, -6173, 5272, 6362, -5045, -6544, 4808, 6716, -4568, -6881, 4319, 7035, -4067, -7183, 3807, 7319, -3544, 
---7448, 3274, 7565, -3002, -7675, 2724, 7772, -2444, -7861, 2159, 7939, -1872, -8007, 1581, 8064, -1290, -8111, 994, 8147, -700, -8173, 402, 8187, -105, -8191, -194, 8183, 490, -8166, -789, 
--8137, 1084, -8098, -1381, 8047, 1673, -7987, -1966, 7914, 2254, -7833, -2542, 7739, 2824, -7636, -3104, 7522, 3379, -7399, -3651, 7264, 3917, -7121, -4179, 6967, 4434, -6805, -4685, 6631, 4928, 
---6451, -5166, 6260, 5396, -6062, -5620, 5854, 5835, -5640, -6044, 5416, 6243, -5186, -6436, 4947, 6618, -4703, -6793, 4451, 6957, -4194, -7113, 3930, 7258, -3661, -7394, 3386, 7519, -3108, -7636, 
--2823, 7740, -2536, -7835, 2244, 7917, -1950, -7991, 1652, 8052, -1352, -8103, 1049, 8141, -746, -8170, 440, 8185, -135, -8191, -172, 8184, 477, -8167, -784, 8137, 1088, -8097, -1392, 8044, 
--1693, -7981, -1994, 7905, 2290, -7820, -2585, 7722, 2874, -7615, -3162, 7495, 3443, -7366, -3722, 7225, 3993, -7075, -4261, 6914, 4521, -6744, -4777, 6562, 5024, -6373, -5266, 6173, 5499, -5966, 
---5726, 5748, 5942, -5524, -6153, 5289, 6353, -5049, -6545, 4800, 6727, -4545, -6900, 4281, 7062, -4014, -7216, 3738, 7358, -3459, -7490, 3172, 7610, -2883, -7721, 2587, 7819, -2289, -7908, 1986, 
--7983, -1682, -8048, 1373, 8099, -1063, -8141, 750, 8169, -438, -8187, 123, 8190, 190, -8184, -506, 8164, 819, -8133, -1133, 8089, 1443, -8034, -1753, 7966, 2059, -7887, -2364, 7795, 2664, 
---7693, -2962, 7578, 3254, -7453, -3543, 7315, 3825, -7168, -4103, 7008, 4374, -6840, -4640, 6659, 4897, -6470, -5149, 6269, 5392, -6061, -5628, 5841, 5854, -5614, -6073, 5377, 6282, -5133, -6483, 
--4880, 6672, -4621, -6853, 4352, 7022, -4079, -7182, 3798, 7329, -3512, -7468, 3219, 7593, -2923, -7708, 2620, 7810, -2316, -7901, 2005, 7979, -1693, -8046, 1376, 8099, -1059, -8142, 738, 8170, 
---418, -8187, 95, 8190, 227, -8182, -550, 8160, 871, -8126, -1192, 8078, 1510, -8020, -1828, 7946, 2141, -7863, -2452, 7765, 2759, -7657, -3063, 7534, 3360, -7402, -3655, 7256, 3941, -7101, 
---4224, 6932, 4498, -6755, -4768, 6564, 5028, -6365, -5282, 6154, 5526, -5935, -5763, 5705, 5989, -5467, -6208, 5218, 6416, -4963, -6615, 4698, 6801, -4427, -6979, 4147, 7144, -3862, -7300, 3569, 
--7442, -3272, -7574, 2968, 7692, -2660, -7799, 2346, 7893, -2030, -7975, 1709, 8043, -1387, -8100, 1060, 8141, -733, -8172, 403, 8187, -74, -8191, -257, 8180, 586, -8157, -916, 8119, 1243, 
---8070, -1570, 8005, 1893, -7930, -2215, 7839, 2531, -7738, -2846, 7621, 3153, -7494, -3458, 7353, 3756, -7202, -4049, 7036, 4334, -6861, -4614, 6672, 4885, -6475, -5149, 6264, 5403, -6045, -5650, 
--5814, 5887, -5574, -6115, 5324, 6331, -5066, -6539, 4798, 6734, -4524, -6920, 4240, 7093, -3950, -7256, 3652, 7404, -3350, -7542, 3040, 7666, -2726, -7779, 2406, 7877, -2083, -7963, 1755, 8035, 
---1426, -8094, 1091, 8138, -757, -8170, 420, 8187, -83, -8191, -255, 8180, 592, -8156, -930, 8117, 1264, -8065, -1599, 7998, 1928, -7920, -2257, 7825, 2580, -7719, -2901, 7598, 3215, -7466, 
---3526, 7318, 3829, -7160, -4127, 6988, 4416, -6805, -4700, 6609, 4974, -6403, -5242, 6184, 5498, -5955, -5748, 5715, 5985, -5466, -6214, 5206, 6430, -4938, -6638, 4660, 6831, -4375, -7015, 4081, 
--7185, -3781, -7344, 3473, 7489, -3160, -7622, 2839, 7740, -2515, -7847, 2185, 7938, -1853, -8017, 1515, 8079, -1176, -8130, 833, 8164, -490, -8185, 144, 8190, 200, -8183, -546, 8159, 889, 
---8122, -1233, 8069, 1573, -8004, -1912, 7922, 2246, -7828, -2578, 7718, 2904, -7596, -3227, 7458, 3542, -7309, -3853, 7145, 4155, -6969, -4452, 6779, 4739, -6579, -5020, 6364, 5289, -6140, -5552, 
--5903, 5802, -5657, -6044, 5398, 6273, -5132, -6493, 4854, 6699, -4569, -6895, 4273, 7077, -3972, -7248, 3661, 7403, -3345, -7547, 3021, 7676, -2693, -7792, 2358, 7892, -2021, -7980, 1678, 8051, 
---1333, -8109, 984, 8150, -635, -8179, 282, 8190, 70, -8188, -423, 8169, 774, -8136, -1125, 8087, 1473, -8024, -1820, 7945, 2162, -7852, -2502, 7743, 2836, -7622, -3167, 7484, 3489, -7334, 
---3808, 7168, 4117, -6990, -4421, 6798, 4715, -6594, -5002, 6376, 5278, -6148, -5546, 5906, 5802, -5655, -6048, 5391, 6282, -5118, -6506, 4834, 6715, -4543, -6914, 4240, 7098, -3932, -7271, 3613, 
--7427, -3290, -7572, 2958, 7700, -2623, -7816, 2280, 7915, -1935, -8000, 1583, 8069, -1231, -8124, 874, 8161, -517, -8185, 157, 8190, 202, -8183, -562, 8157, 920, -8117, -1278, 8060, 1631, 
---7989, -1984, 7901, 2331, -7799, -2676, 7680, 3013, -7549, -3347, 7400, 3673, -7239, -3994, 7061, 4305, -6872, -4610, 6667, 4904, -6451, -5190, 6220, 5465, -5979, -5731, 5724, 5983, -5460, -6227, 
--5183, 6456, -4897, -6674, 4599, 6877, -4295, -7069, 3979, 7245, -3658, -7409, 3327, 7556, -2992, -7691, 2648, 7808, -2301, -7911, 1947, 7997, -1591, -8069, 1230, 8123, -868, -8163, 502, 8184, 
---137, -8191, -231, 8180, 596, -8154, -963, 8110, 1325, -8052, -1687, 7975, 2044, -7884, -2399, 7776, 2747, -7653, -3092, 7513, 3429, -7360, -3761, 7190, 4084, -7007, -4401, 6807, 4707, -6596, 
---5005, 6369, 5291, -6132, -5569, 5879, 5834, -5617, -6088, 5340, 6329, -5055, -6559, 4757, 6773, -4452, -6976, 4135, 7162, -3811, -7336, 3478, 7492, -3139, -7636, 2791, 7762, -2439, -7873, 2081, 
--7967, -1719, -8046, 1352, 8107, -985, -8152, 612, 8179, -241, -8191, -134, 8184, 506, -8162, -880, 8121, 1249, -8065, -1619, 7990, 1983, -7900, -2345, 7792, 2701, -7669, -3053, 7529, 3397, 
---7374, -3736, 7202, 4065, -7016, -4388, 6814, 4699, -6599, -5003, 6368, 5295, -6126, -5578, 5869, 5847, -5601, -6105, 5319, 6349, -5027, -6582, 4723, 6798, -4410, -7003, 4086, 7190, -3756, -7365, 
--3415, 7522, -3068, -7664, 2713, 7789, -2354, -7899, 1987, 7990, -1618, -8065, 1244, 8122, -868, -8163, 489, 8185, -110, -8191, -271, 8178, 650, -8148, -1030, 8099, 1405, -8035, -1780, 7951, 
--2149, -7852, -2515, 7734, 2875, -7601, -3230, 7450, 3576, -7284, -3917, 7100, 4248, -6903, -4571, 6688, 4883, -6461, -5186, 6217, 5475, -5962, -5755, 5692, 6021, -5411, -6275, 5116, 6514, -4811, 
---6741, 4494, 6951, -4169, -7147, 3832, 7326, -3489, -7491, 3136, 7638, -2778, -7770, 2411, 7882, -2041, -7979, 1664, 8057, -1286, -8118, 902, 8160, -518, -8185, 131, 8190, 255, -8179, -643, 
--8148, 1027, -8100, -1411, 8033, 1790, -7949, -2167, 7845, 2538, -7726, -2905, 7587, 3264, -7433, -3617, 7261, 3961, -7074, -4298, 6869, 4623, -6650, -4940, 6414, 5244, -6166, -5539, 5901, 5819, 
---5625, -6087, 5334, 6341, -5033, -6582, 4718, 6806, -4394, -7016, 4058, 7209, -3715, -7388, 3361, 7547, -3001, -7692, 2632, 7817, -2259, -7926, 1878, 8015, -1495, -8087, 1107, 8140, -717, -8175, 
--324, 8189, 68, -8187, -462, 8164, 853, -8124, -1245, 8063, 1632, -7986, -2017, 7888, 2396, -7773, -2771, 7639, 3138, -7488, -3500, 7319, 3853, -7134, -4198, 6930, 4532, -6712, -4857, 6476, 
--5169, -6227, -5471, 5962, 5759, -5684, -6035, 5391, 6295, -5087, -6542, 4769, 6773, -4441, -6989, 4101, 7187, -3753, -7370, 3394, 7534, -3029, -7682, 2655, 7810, -2276, -7922, 1889, 8013, -1500, 
---8087, 1105, 8140, -709, -8176, 310, 8190, 89, -8186, -489, 8162, 887, -8119, -1285, 8055, 1677, -7974, -2068, 7872, 2453, -7753, -2833, 7613, 3205, -7457, -3571, 7281, 3927, -7090, -4276, 
--6879, 4613, -6654, -4940, 6410, 5254, -6153, -5558, 5879, 5846, -5592, -6122, 5290, 6381, -4977, -6627, 4649, 6855, -4313, -7069, 3963, 7263, -3606, -7442, 3238, 7601, -2863, -7743, 2480, 7865, 
---2092, -7969, 1697, 8052, -1300, -8117, 897, 8161, -494, -8186, 87, 8190, 318, -8175, -724, 8138, 1127, -8083, -1529, 8006, 1926, -7911, -2320, 7795, 2706, -7662, -3088, 7507, 3461, -7336, 
---3827, 7144, 4182, -6937, -4529, 6710, 4862, -6469, -5186, 6209, 5495, -5936, -5792, 5645, 6073, -5343, -6341, 5025, 6591, -4696, -6827, 4354, 7044, -4002, -7245, 3638, 7427, -3267, -7591, 2886, 
--7735, -2499, -7862, 2103, 7966, -1704, -8053, 1299, 8117, -892, -8163, 480, 8186, -70, -8190, -344, 8172, 754, -8135, -1165, 8075, 1571, -7997, -1975, 7897, 2372, -7778, -2766, 7637, 3150, 
---7479, -3529, 7300, 3897, -7104, -4257, 6888, 4605, -6655, -4943, 6404, 5266, -6139, -5578, 5855, 5874, -5558, -6157, 5245, 6422, -4920, -6672, 4580, 6904, -4231, -7120, 3868, 7316, -3497, -7494, 
--3115, 7652, -2726, -7792, 2329, 7909, -1927, -8008, 1518, 8085, -1106, -8142, 690, 8176, -274, -8191, -146, 8183, 563, -8155, -980, 8104, 1394, -8034, -1806, 7940, 2211, -7828, -2613, 7693, 
--3006, -7540, -3393, 7365, 3770, -7173, -4139, 6960, 4495, -6730, -4842, 6480, 5174, -6215, -5494, 5932, 5798, -5635, -6089, 5320, 6362, -4994, -6620, 4652, 6859, -4300, -7081, 3934, 7283, -3559, 
---7468, 3173, 7630, -2780, -7775, 2377, 7897, -1970, -7999, 1556, 8079, -1139, -8139, 717, 8175, -294, -8191, -131, 8183, 554, -8156, -978, 8104, 1397, -8032, -1815, 7937, 2226, -7823, -2633, 
--7685, 3031, -7528, -3424, 7349, 3805, -7152, -4178, 6934, 4538, -6699, -4888, 6443, 5223, -6172, -5545, 5882, 5851, -5578, -6143, 5256, 6416, -4922, -6674, 4572, 6912, -4212, -7134, 3838, 7333, 
---3456, -7515, 3061, 7674, -2660, -7815, 2250, 7931, -1835, -8029, 1414, 8102, -990, -8155, 561, 8183, -132, -8191, -299, 8174, 728, -8137, -1157, 8075, 1580, -7993, -2002, 7887, 2416, -7761, 
---2826, 7611, 3226, -7442, -3619, 7250, 4001, -7040, -4373, 6808, 4731, -6559, -5079, 6290, 5410, -6005, -5729, 5701, 6029, -5383, -6315, 5048, 6581, -4700, -6831, 4338, 7060, -3964, -7271, 3578, 
--7460, -3183, -7630, 2777, 7776, -2366, -7903, 1945, 8005, -1520, -8087, 1090, 8144, -657, -8180, 221, 8190, 214, -8180, -650, 8144, 1083, -8088, -1516, 8006, 1942, -7903, -2364, 7776, 2778, 
---7629, -3187, 7458, 3584, -7267, -3974, 7054, 4350, -6822, -4716, 6569, 5066, -6298, -5405, 6008, 5725, -5702, -6032, 5378, 6319, -5040, -6591, 4685, 6841, -4319, -7074, 3938, 7285, -3548, -7476, 
--3145, 7644, -2735, -7792, 2315, 7916, -1889, -8019, 1457, 8096, -1021, -8152, 581, 8183, -141, -8191, -302, 8174, 742, -8135, -1182, 8070, 1617, -7984, -2050, 7872, 2474, -7739, -2894, 7581, 
--3303, -7404, -3705, 7202, 4094, -6981, -4473, 6738, 4837, -6476, -5190, 6194, 5525, -5895, -5846, 5577, 6148, -5244, -6433, 4893, 6698, -4530, -6946, 4151, 7171, -3762, -7376, 3360, 7558, -2949, 
---7720, 2527, 7857, -2100, -7972, 1664, 8062, -1225, -8130, 781, 8171, -336, -8191, -113, 8184, 559, -8154, -1006, 8098, 1448, -8020, -1888, 7915, 2320, -7789, -2748, 7638, 3165, -7465, -3576, 
--7268, 3973, -7051, -4361, 6811, 4734, -6552, -5095, 6271, 5439, -5973, -5768, 5655, 6078, -5322, -6372, 4970, 6644, -4605, -6899, 4225, 7130, -3833, -7343, 3427, 7531, -3013, -7698, 2587, 7840, 
---2155, -7959, 1715, 8053, -1271, -8124, 821, 8169, -370, -8190, -84, 8185, 536, -8156, -988, 8100, 1436, -8022, -1881, 7916, 2319, -7789, -2752, 7635, 3175, -7460, -3590, 7260, 3992, -7039, 
---4384, 6794, 4761, -6531, -5125, 6245, 5471, -5941, -5803, 5617, 6115, -5278, -6410, 4920, 6683, -4548, -6937, 4160, 7168, -3761, -7379, 3349, 7565, -2927, -7730, 2494, 7868, -2056, -7984, 1608, 
--8073, -1158, -8139, 702, 8177, -245, -8191, -215, 8178, 672, -8142, -1129, 8077, 1581, -7990, -2031, 7875, 2472, -7737, -2907, 7573, 3331, -7387, -3747, 7175, 4150, -6943, -4541, 6686, 4916, 
---6411, -5278, 6112, 5621, -5797, -5949, 5461, 6256, -5109, -6545, 4739, 6811, -4355, -7058, 3956, 7280, -3546, -7482, 3122, 7657, -2691, -7810, 2248, 7936, -1800, -8039, 1344, 8114, -886, -8165, 
--422, 8188, 41, -8187, -506, 8157, 967, -8103, -1428, 8021, 1882, -7915, -2333, 7782, 2774, -7625, -3208, 7442, 3630, -7237, -4043, 7006, 4441, -6754, -4826, 6478, 5194, -6183, -5547, 5866, 
--5881, -5532, -6197, 5177, 6491, -4808, -6767, 4421, 7018, -4021, -7249, 3606, 7454, -3181, -7637, 2743, 7793, -2298, -7925, 1844, 8030, -1385, -8110, 920, 8162, -453, -8189, -18, 8187, 486, 
---8160, -955, 8104, 1419, -8023, -1881, 7914, 2335, -7781, -2783, 7620, 3220, -7436, -3649, 7225, 4063, -6992, -4467, 6734, 4854, -6456, -5227, 6154, 5580, -5833, -5918, 5491, 6233, -5132, -6530, 
--4754, 6804, -4362, -7057, 3953, 7284, -3533, -7489, 3099, 7668, -2657, -7822, 2203, 7949, -1744, -8051, 1277, 8124, -807, -8172, 333, 8190, 141, -8183, -617, 8146, 1089, -8084, -1559, 7992, 
--2022, -7876, -2481, 7731, 2929, -7561, -3370, 7364, 3797, -7144, -4214, 6898, 4615, -6630, -5002, 6338, 5370, -6026, -5723, 5691, 6054, -5339, -6366, 4966, 6655, -4579, -6923, 4174, 7166, -3756, 
---7387, 3323, 7580, -2881, -7749, 2426, 7890, -1966, -8006, 1496, 8093, -1023, -8154, 544, 8185, -65, -8190, -416, 8164, 894, -8113, -1371, 8031, 1842, -7924, -2308, 7787, 2765, -7626, -3214, 
--7436, 3651, -7222, -4077, 6981, 4487, -6718, -4883, 6430, 5261, -6121, -5623, 5788, 5963, -5437, -6285, 5066, 6582, -4678, -6860, 4272, 7111, -3853, -7340, 3418, 7541, -2974, -7717, 2516, 7865, 
---2052, -7988, 1578, 8080, -1101, -8146, 617, 8182, -133, -8191, -353, 8169, 837, -8120, -1319, 8041, 1796, -7935, -2268, 7800, 2730, -7638, -3185, 7448, 3627, -7233, -4058, 6991, 4473, -6726, 
---4875, 6435, 5257, -6122, -5622, 5786, 5966, -5432, -6291, 5056, 6592, -4663, -6871, 4252, 7124, -3828, -7353, 3388, 7555, -2937, -7731, 2474, 7878, -2004, -7999, 1525, 8089, -1041, -8153, 552, 
--8185, -63, -8189, -429, 8163, 917, -8109, -1404, 8024, 1885, -7911, -2360, 7769, 2826, -7600, -3283, 7402, 3727, -7179, -4160, 6928, 4575, -6654, -4977, 6353, 5358, -6032, -5722, 5686, 6064, 
---5322, -6385, 4936, 6682, -4534, -6956, 4113, 7203, -3680, -7426, 3230, 7620, -2771, -7789, 2300, 7927, -1822, -8038, 1335, 8118, -845, -8170, 349, 8190, 146, -8182, -642, 8142, 1134, -8074, 
---1625, 7975, 2107, -7848, -2584, 7690, 3050, -7506, -3507, 7292, 3948, -7054, -4378, 6787, 4789, -6496, -5185, 6180, 5560, -5843, -5917, 5482, 6249, -5102, -6561, 4702, 6847, -4285, -7109, 3851, 
--7342, -3404, -7551, 2943, 7730, -2472, -7882, 1990, 8002, -1502, -8095, 1007, 8155, -509, -8187, 7, 8187, 492, -8158, -993, 8096, 1487, -8006, -1978, 7884, 2461, -7734, -2936, 7553, 3398, 
---7346, -3849, 7108, 4284, -6846, -4706, 6557, 5107, -6244, -5492, 5905, 5854, -5547, -6196, 5165, 6513, -4765, -6807, 4345, 7073, -3910, -7315, 3459, 7527, -2996, -7713, 2520, 7867, -2036, -7994, 
--1541, 8088, -1043, -8153, 539, 8185, -34, -8189, -473, 8158, 976, -8099, -1478, 8007, 1972, -7886, -2461, 7732, 2938, -7551, -3407, 7339, 3861, -7101, -4302, 6833, 4725, -6541, -5131, 6222, 
--5516, -5881, -5882, 5515, 6224, -5129, -6544, 4721, 6836, -4298, -7104, 3855, 7343, -3399, -7555, 2928, 7737, -2447, -7890, 1955, 8011, -1457, -8102, 951, 8161, -443, -8189, -69, 8184, 579, 
---8149, -1088, 8080, 1592, -7982, -2091, 7850, 2581, -7690, -3063, 7497, 3531, -7277, -3987, 7027, 4426, -6751, -4849, 6446, 5252, -6118, -5637, 5764, 5997, -5389, -6336, 4990, 6648, -4574, -6936, 
--4138, 7195, -3687, -7427, 3219, 7629, -2741, -7802, 2250, 7942, -1751, -8053, 1243, 8131, -733, -8178, 217, 8190, 298, -8173, -814, 8120, 1325, -8038, -1833, 7921, 2332, -7775, -2823, 7596, 
--3302, -7388, -3769, 7149, 4220, -6884, -4656, 6588, 5072, -6268, -5469, 5922, 5843, -5553, -6195, 5160, 6521, -4747, -6823, 4314, 7095, -3865, -7341, 3399, 7556, -2921, -7742, 2428, 7895, -1928, 
---8019, 1418, 8108, -904, -8166, 384, 8190, 136, -8182, -657, 8139, 1174, -8065, -1688, 7957, 2194, -7818, -2693, 7646, 3179, -7444, -3655, 7210, 4113, -6949, -4558, 6657, 4982, -6340, -5387, 
--5995, 5769, -5627, -6130, 5235, 6463, -4823, -6773, 4388, 7052, -3938, -7305, 3470, 7526, -2989, -7719, 2494, 7877, -1990, -8006, 1476, 8100, -957, -8162, 433, 8189, 92, -8184, -618, 8143, 
--1140, -8071, -1659, 7963, 2170, -7825, -2674, 7652, 3165, -7449, -3645, 7214, 4109, -6950, -4557, 6656, 4985, -6336, -5394, 5987, 5779, -5616, -6142, 5219, 6478, -4802, -6788, 4363, 7069, -3907, 
---7322, 3433, 7543, -2947, -7734, 2446, 7892, -1937, -8018, 1417, 8109, -893, -8167, 364, 8190, 166, -8180, -697, 8134, 1223, -8056, -1746, 7942, 2260, -7796, -2767, 7615, 3260, -7405, -3742, 
--7161, 4206, -6889, -4654, 6585, 5081, -6256, -5489, 5898, 5872, -5517, -6232, 5110, 6563, -4684, -6869, 4236, 7144, -3771, -7391, 3289, 7604, -2794, -7787, 2285, 7936, -1768, -8052, 1242, 8132, 
---712, -8179, 176, 8190, 358, -8168, -893, 8108, 1422, -8016, -1947, 7888, 2463, -7728, -2969, 7532, 3462, -7306, -3941, 7047, 4402, -6760, -4846, 6441, 5268, -6096, -5669, 5723, 6043, -5328, 
---6394, 4907, 6715, -4466, -7010, 4005, 7272, -3528, -7505, 3033, 7704, -2527, -7871, 2008, 8002, -1482, -8101, 948, 8162, -411, -8190, -130, 8181, 668, -8138, -1206, 8057, 1736, -7944, -2262, 
--7793, 2775, -7611, -3279, 7393, 3767, -7145, -4240, 6864, 4693, -6555, -5127, 6215, 5538, -5849, -5926, 5456, 6286, -5040, -6621, 4601, 6925, -4143, -7200, 3664, 7442, -3172, -7654, 2663, 7830, 
---2144, -7973, 1614, 8079, -1078, -8152, 535, 8186, 8, -8187, -553, 8149, 1094, -8077, -1633, 7967, 2162, -7824, -2684, 7645, 3193, -7433, -3689, 7186, 4167, -6909, -4629, 6599, 5068, -6262, 
---5487, 5895, 5880, -5503, -6248, 5085, 6587, -4646, -6898, 4184, 7177, -3705, -7426, 3207, 7639, -2697, -7821, 2172, 7965, -1640, -8076, 1098, 8149, -553, -8187, 3, 8186, 545, -8150, -1093, 
--8076, 1634, -7967, -2170, 7821, 2694, -7641, -3208, 7424, 3706, -7176, -4190, 6893, 4652, -6581, -5096, 6237, 5515, -5867, -5911, 5468, 6278, -5046, -6619, 4599, 6928, -4133, -7208, 3646, 7453, 
---3144, -7666, 2626, 7842, -2097, -7985, 1557, 8089, -1012, -8158, 459, 8188, 93, -8183, -648, 8138, 1197, -8058, -1744, 7939, 2280, -7786, -2808, 7595, 3322, -7371, -3822, 7110, 4304, -6820, 
---4767, 6495, 5207, -6143, -5625, 5760, 6015, -5353, -6379, 4918, 6712, -4463, -7017, 3985, 7287, -3491, -7525, 2978, 7727, -2453, -7895, 1915, 8024, -1369, -8118, 815, 8173, -259, -8191, -300, 
--8170, 856, -8113, -1411, 8015, 1957, -7883, -2496, 7711, 3021, -7506, -3535, 7264, 4031, -6989, -4509, 6680, 4965, -6341, -5400, 5971, 5808, -5574, -6190, 5149, 6542, -4702, -6865, 4231, 7154, 
---3741, -7411, 3232, 7632, -2710, -7819, 2172, 7967, -1626, -8080, 1071, 8152, -512, -8188, -52, 8184, 613, -8143, -1174, 8061, 1728, -7943, -2275, 7785, 2810, -7593, -3334, 7362, 3840, -7099, 
---4330, 6799, 4798, -6470, -5245, 6107, 5665, -5717, -6061, 5298, 6425, -4855, -6761, 4387, 7064, -3900, -7334, 3393, 7567, -2870, -7767, 2332, 7927, -1785, -8052, 1227, 8136, -664, -8183, 97, 
--8188, 469, -8157, -1036, 8084, 1595, -7974, -2149, 7824, 2691, -7639, -3222, 7414, 3736, -7156, -4234, 6861, 4709, -6534, -5164, 6174, 5593, -5787, -5996, 5369, 6368, -4926, -6712, 4458, 7022, 
---3970, -7299, 3461, 7539, -2937, -7745, 2396, 7911, -1845, -8040, 1284, 8129, -718, -8180, 146, 8189, 425, -8161, -996, 8090, 1560, -7982, -2119, 7833, 2666, -7647, -3202, 7423, 3720, -7163, 
---4222, 6867, 4702, -6538, -5161, 6176, 5593, -5785, -5999, 5364, 6374, -4918, -6720, 4445, 7031, -3953, -7309, 3439, 7550, -2910, -7755, 2364, 7920, -1809, -8048, 1242, 8134, -671, -8183, 95, 
--8188, 480, -8155, -1055, 8080, 1623, -7967, -2185, 7812, 2735, -7620, -3273, 7388, 3793, -7122, -4296, 6818, 4776, -6482, -5234, 6111, 5665, -5712, -6069, 5283, 6442, -4829, -6784, 4348, 7090, 
---3848, -7363, 3326, 7598, -2789, -7796, 2237, 7953, -1674, -8073, 1102, 8150, -525, -8188, -56, 8183, 635, -8139, -1213, 8052, 1784, -7926, -2347, 7759, 2897, -7554, -3435, 7309, 3953, -7029, 
---4453, 6712, 4930, -6362, -5383, 5978, 5807, -5566, -6204, 5124, 6568, -4657, -6901, 4164, 7196, -3653, -7458, 3120, 7679, -2574, -7864, 2012, 8006, -1442, -8110, 862, 8171, -280, -8191, -306, 
--8169, 889, -8106, -1469, 8000, 2040, -7855, -2603, 7668, 3151, -7444, -3684, 7179, 4197, -6879, -4691, 6542, 5158, -6174, -5602, 5771, 6014, -5341, -6398, 4881, 6748, -4398, -7064, 3890, 7342, 
---3364, -7585, 2819, 7786, -2260, -7950, 1688, 8070, -1109, -8151, 522, 8187, 66, -8184, -656, 8135, 1241, -8047, -1821, 7915, 2390, -7744, -2949, 7530, 3491, -7279, -4017, 6989, 4520, -6664, 
---5002, 6302, 5455, -5909, -5883, 5483, 6278, -5031, -6642, 4550, 6970, -4047, -7264, 3521, 7518, -2978, -7734, 2417, 7908, -1846, -8042, 1263, 8133, -675, -8183, 81, 8188, 512, -8152, -1103, 
--8071, 1688, -7949, -2265, 7784, 2829, -7579, -3381, 7333, 3912, -7050, -4425, 6727, 4913, -6371, -5377, 5979, 5811, -5558, -6216, 5104, 6587, -4626, -6924, 4121, 7223, -3596, -7486, 3050, 7707, 
---2489, -7890, 1913, 8028, -1328, -8126, 735, 8179, -139, -8190, -460, 8155, 1054, -8079, -1645, 7958, 2226, -7797, -2797, 7591, 3351, -7347, -3889, 7062, 4405, -6740, -4899, 6381, 5365, -5989, 
---5805, 5563, 6211, -5109, -6586, 4625, 6924, -4118, -7227, 3587, 7490, -3039, -7714, 2472, 7894, -1893, -8034, 1302, 8129, -706, -8181, 104, 8188, 497, -8153, -1097, 8071, 1690, -7948, -2276, 
--7779, 2848, -7570, -3406, 7319, 3944, -7029, -4463, 6699, 4956, -6335, -5424, 5934, 5860, -5503, -6267, 5039, 6638, -4550, -6975, 4034, 7272, -3498, -7531, 2941, 7748, -2369, -7924, 1783, 8055, 
---1188, -8143, 585, 8186, 20, -8185, -627, 8138, 1229, -8048, -1826, 7911, 2411, -7734, -2985, 7511, 3541, -7250, -4080, 6946, 4594, -6606, -5086, 6228, 5547, -5817, -5980, 5372, 6378, -4899, 
---6743, 4397, 7069, -3872, -7358, 3324, 7604, -2759, -7810, 2177, 7971, -1584, -8090, 981, 8162, -374, -8191, -237, 8173, 846, -8110, -1451, 8001, 2047, -7849, -2634, 7652, 3204, -7414, -3759, 
--7132, 4290, -6813, -4800, 6453, 5281, -6059, -5735, 5629, 6155, -5170, -6543, 4679, 6892, -4165, -7205, 3624, 7475, -3065, -7706, 2487, 7891, -1897, -8034, 1293, 8130, -685, -8183, 70, 8187, 
--543, -8147, -1156, 8060, 1760, -7928, -2357, 7750, 2938, -7531, -3505, 7266, 4050, -6963, -4575, 6617, 5071, -6237, -5542, 5819, 5979, -5370, -6384, 4888, 6751, -4380, -7082, 3846, 7371, -3291, 
---7620, 2715, 7824, -2126, -7985, 1523, 8099, -912, -8169, 294, 8190, 323, -8167, -941, 8095, 1552, -7979, -2156, 7815, 2746, -7608, -3323, 7355, 3878, -7063, -4414, 6728, 4922, -6356, -5405, 
--5946, 5854, -5503, -6272, 5026, 6652, -4523, -6996, 3991, 7298, -3439, -7560, 2864, 7777, -2274, -7950, 1670, 8076, -1057, -8157, 436, 8190, 186, -8176, -808, 8114, 1425, -8007, -2035, 7851, 
--2631, -7651, -3215, 7406, 3778, -7119, -4321, 6788, 4838, -6421, -5328, 6013, 5786, -5573, -6212, 5098, 6600, -4595, -6952, 4064, 7261, -3510, -7530, 2934, 7753, -2342, -7933, 1735, 8065, -1119, 
---8152, 495, 8188, 131, -8179, -758, 8120, 1378, -8016, -1993, 7862, 2595, -7664, -3183, 7419, 3751, -7133, -4299, 6802, 4819, -6433, -5314, 6025, 5776, -5582, -6205, 5105, 6596, -4599, -6950, 
--4064, 7262, -3507, -7532, 2927, 7756, -2331, -7937, 1720, 8068, -1100, -8154, 471, 8189, 159, -8178, -790, 8116, 1414, -8008, -2032, 7850, 2636, -7648, -3227, 7398, 3797, -7106, -4346, 6770, 
--4868, -6395, -5363, 5980, 5824, -5531, -6252, 5046, 6641, -4534, -6993, 3992, 7301, -3428, -7567, 2842, 7786, -2240, -7960, 1623, 8085, -998, -8163, 364, 8190, 269, -8170, -904, 8099, 1531, 
---7982, -2151, 7814, 2756, -7601, -3347, 7340, 3916, -7037, -4464, 6689, 4982, -6303, -5473, 5877, 5929, -5417, -6351, 4922, 6733, -4399, -7076, 3847, 7375, -3274, -7631, 2679, 7838, -2069, -8001, 
--1445, 8112, -813, -8177, 175, 8189, 463, -8154, -1100, 8067, 1728, -7933, -2349, 7749, 2953, -7519, -3541, 7242, 4106, -6922, -4648, 6558, 5160, -6155, -5642, 5713, 6088, -5237, -6499, 4728, 
--6868, -4191, -7197, 3626, 7480, -3041, -7719, 2435, 7909, -1816, -8053, 1184, 8145, -546, -8188, -97, 8180, 738, -8123, -1377, 8014, 2005, -7857, -2624, 7650, 3224, -7398, -3806, 7097, 4363, 
---6755, -4896, 6369, 5396, -5946, -5865, 5483, 6295, -4988, -6689, 4460, 7040, -3907, -7348, 3327, 7610, -2728, -7826, 2110, 7991, -1480, -8109, 840, 8174, -195, -8190, -452, 8154, 1095, -8068, 
---1734, 7930, 2359, -7745, -2973, 7509, 3565, -7228, -4138, 6899, 4683, -6530, -5201, 6117, 5684, -5668, -6134, 5181, 6543, -4664, -6914, 4115, 7239, -3542, -7521, 2945, 7754, -2330, -7939, 1699, 
--8073, -1060, -8158, 411, 8190, 239, -8172, -889, 8100, 1532, -7980, -2167, 7806, 2787, -7586, -3391, 7315, 3972, -7000, -4530, 6638, 5058, -6237, -5555, 5793, 6016, -5315, -6440, 4800, 6822, 
---4258, -7163, 3685, 7456, -3092, -7703, 2476, 7900, -1846, -8048, 1203, 8143, -553, -8188, -102, 8179, 754, -8120, -1404, 8007, 2044, -7844, -2672, 7629, 3282, -7368, -3872, 7057, 4436, -6703, 
---4974, 6303, 5478, -5865, -5949, 5388, 6380, -4877, -6772, 4333, 7118, -3763, -7421, 3167, 7674, -2552, -7880, 1918, 8033, -1274, -8137, 619, 8185, 38, -8183, -696, 8126, 1349, -8019, -1995, 
--7857, 2626, -7647, -3242, 7385, 3836, -7077, -4407, 6721, 4947, -6324, -5458, 5883, 5931, -5406, -6368, 4891, 6761, -4347, -7113, 3772, 7416, -3174, -7674, 2554, 7879, -1919, -8035, 1269, 8136, 
---612, -8187, -51, 8182, 711, -8125, -1369, 8013, 2017, -7851, -2653, 7635, 3270, -7372, -3868, 7057, 4439, -6699, -4982, 6294, 5491, -5850, -5967, 5365, 6401, -4847, -6795, 4295, 7142, -3716, 
---7445, 3111, 7697, -2487, -7900, 1844, 8048, -1191, -8146, 528, 8188, 136, -8178, -802, 8112, 1461, -7994, -2113, 7821, 2748, -7598, -3368, 7323, 3963, -7001, -4535, 6631, 5074, -6218, -5582, 
--5762, 6051, -5270, -6482, 4740, 6867, -4180, -7209, 3591, 7502, -2980, -7746, 2346, 7937, -1699, -8076, 1038, 8160, -372, -8191, -299, 8166, 966, -8088, -1629, 7954, 2279, -7768, -2916, 7528, 
--3531, -7240, -4125, 6901, 4690, -6518, -5225, 6089, 5723, -5620, -6185, 5112, 6603, -4571, -6979, 3998, 7307, -3399, -7587, 2775, 7813, -2134, -7990, 1477, 8110, -811, -8178, 138, 8188, 535, 
---8145, -1206, 8045, 1867, -7892, -2517, 7684, 3149, -7426, -3761, 7115, 4347, -6758, -4904, 6353, 5427, -5906, -5915, 5417, 6361, -4894, -6766, 4335, 7122, -3748, -7433, 3133, 7690, -2499, -7898, 
--1846, 8049, -1181, -8148, 507, 8189, 169, -8176, -846, 8105, 1516, -7980, -2177, 7799, 2822, -7567, -3449, 7280, 4051, -6945, -4628, 6561, 5170, -6133, -5680, 5661, 6148, -5153, -6577, 4606, 
--6958, -4030, -7293, 3423, 7576, -2795, -7809, 2146, 7987, -1483, -8111, 808, 8177, -129, -8189, -552, 8142, 1229, -8041, -1899, 7882, 2554, -7670, -3193, 7403, 3809, -7087, -4400, 6720, 4959, 
---6307, -5485, 5849, 5972, -5352, -6419, 4816, 6820, -4248, -7175, 3648, 7479, -3025, -7732, 2378, 7930, -1717, -8074, 1041, 8160, -360, -8191, -325, 8163, 1007, -8080, -1684, 7938, 2347, -7743, 
---2996, 7491, 3622, -7189, -4225, 6834, 4797, -6433, -5336, 5985, 5837, -5497, -6299, 4968, 6714, -4405, -7085, 3810, 7404, -3190, -7672, 2545, 7885, -1884, -8044, 1207, 8145, -524, -8190, -166, 
--8175, 852, -8104, -1534, 7974, 2204, -7790, -2860, 7548, 3495, -7255, -4106, 6908, 4687, -6514, -5237, 6072, 5747, -5589, -6219, 5064, 6645, -4504, -7026, 3911, 7355, -3291, -7634, 2646, 7856, 
---1984, -8024, 1306, 8134, -620, -8187, -73, 8180, 763, -8116, -1450, 7993, 2125, -7814, -2787, 7577, 3427, -7288, -4045, 6945, 4632, -6554, -5188, 6113, 5705, -5631, -6183, 5106, 6614, -4546, 
---7001, 3952, 7335, -3331, -7618, 2684, 7845, -2019, -8017, 1337, 8130, -648, -8186, -48, 8181, 742, -8119, -1433, 7996, 2112, -7818, -2777, 7580, 3421, -7290, -4042, 6946, 4632, -6552, -5191, 
--6109, 5710, -5624, -6190, 5096, 6623, -4532, -7010, 3934, 7345, -3309, -7628, 2657, 7854, -1988, -8024, 1303, 8134, -609, -8187, -90, 8179, 788, -8112, -1482, 7985, 2163, -7801, -2831, 7558, 
--3476, -7262, -4098, 6910, 4688, -6510, -5246, 6060, 5764, -5568, -6241, 5032, 6671, -4462, -7055, 3857, 7384, -3225, -7661, 2567, 7881, -1892, -8044, 1201, 8146, -503, -8190, -200, 8172, 901, 
---8096, -1597, 7957, 2279, -7763, -2947, 7508, 3592, -7201, -4212, 6838, 4799, -6426, -5352, 5965, 5864, -5461, -6335, 4915, 6757, -4334, -7131, 3719, 7451, -3078, -7717, 2412, 7924, -1730, -8074, 
--1033, 8162, -330, -8191, -378, 8158, 1080, -8066, -1778, 7911, 2460, -7700, -3126, 7429, 3766, -7104, -4381, 6725, 4961, -6297, -5507, 5820, 6009, -5301, -6469, 4741, 6878, -4146, -7238, 3519, 
--7541, -2867, -7791, 2191, 7979, -1501, -8110, 797, 8178, -89, -8187, -622, 8132, 1326, -8018, -2023, 7842, 2702, -7608, -3364, 7315, 3998, -6969, -4604, 6568, 5174, -6119, -5706, 5623, 6194, 
---5085, -6637, 4507, 7028, -3897, -7368, 3254, 7651, -2590, -7877, 1903, 8042, -1204, -8147, 493, 8189, 220, -8171, -933, 8089, 1637, -7947, -2331, 7743, 3005, -7482, -3659, 7161, 4283, -6789, 
---4877, 6362, 5431, -5889, -5946, 5368, 6414, -4809, -6836, 4210, 7203, -3581, -7517, 2923, 7772, -2244, -7969, 1546, 8103, -838, -8177, 121, 8187, 595, -8136, -1309, 8020, 2011, -7845, -2699, 
--7608, 3365, -7313, -4007, 6961, 4617, -6557, -5193, 6100, 5728, -5598, -6220, 5051, 6663, -4467, -7056, 3846, 7393, -3198, -7675, 2522, 7896, -1829, -8058, 1119, 8155, -403, -8191, -319, 8162, 
--1036, -8072, -1748, 7917, 2444, -7703, -3124, 7427, 3777, -7095, -4403, 6706, 4994, -6266, -5547, 5776, 6056, -5243, -6519, 4667, 6930, -4056, -7289, 3411, 7590, -2742, -7833, 2049, 8013, -1342, 
---8132, 622, 8186, 101, -8178, -825, 8104, 1541, -7969, -2247, 7769, 2934, -7511, -3600, 7191, 4235, -6817, -4840, 6387, 5405, -5909, -5930, 5382, 6406, -4815, -6834, 4208, 7206, -3570, -7524, 
--2901, 7780, -2212, -7978, 1502, 8110, -783, -8181, 55, 8185, 671, -8126, -1394, 8001, 2105, -7815, -2801, 7565, 3472, -7257, -4119, 6889, 4731, -6469, -5308, 5996, 5841, -5476, -6330, 4911, 
--6767, -4309, -7152, 3671, 7478, -3005, -7747, 2313, 7952, -1605, -8096, 882, 8174, -153, -8189, -579, 8136, 1305, -8020, -2022, 7839, 2722, -7597, -3401, 7292, 4052, -6930, -4673, 6511, 5254, 
---6042, -5796, 5523, 6289, -4961, -6734, 4357, 7124, -3720, -7458, 3051, 7730, -2359, -7942, 1646, 8089, -922, -8173, 188, 8189, 545, -8141, -1277, 8025, 1996, -7847, -2701, 7603, 3383, -7300, 
---4040, 6937, 4662, -6519, -5249, 6046, 5791, -5526, -6289, 4960, 6734, -4355, -7127, 3713, 7460, -3042, -7735, 2345, 7945, -1630, -8093, 901, 8173, -165, -8189, -574, 8136, 1306, -8019, -2030, 
--7835, 2736, -7590, -3422, 7280, 4078, -6913, -4703, 6487, 5287, -6011, -5831, 5483, 6326, -4913, -6770, 4300, 7158, -3654, -7489, 2976, 7758, -2275, -7964, 1553, 8104, -821, -8179, 80, 8185, 
--660, -8126, -1397, 7999, 2121, -7808, -2829, 7550, 3513, -7233, -4170, 6854, 4790, -6420, -5373, 5932, 5911, -5397, -6401, 4815, 6838, -4195, -7219, 3538, 7540, -2854, -7800, 2144, 7994, -1419, 
---8124, 679, 8185, 64, -8180, -809, 8105, 1546, -7966, -2272, 7758, 2977, -7488, -3660, 7154, 4310, -6762, -4927, 6312, 5501, -5812, -6032, 5261, 6511, -4668, -6937, 4034, 7305, -3369, -7613, 
--2673, 7856, -1957, -8035, 1222, 8146, -479, -8191, -270, 8165, 1015, -8073, -1754, 7912, 2477, -7686, -3181, 7395, 3856, -7043, -4502, 6630, 5107, -6163, -5673, 5643, 6188, -5077, -6654, 4467, 
--7063, -3820, -7414, 3140, 7701, -2435, -7925, 1707, 8080, -967, -8170, 216, 8189, 534, -8141, -1283, 8022, 2018, -7838, -2739, 7585, 3435, -7270, -4104, 6892, 4737, -6458, -5332, 5966, 5879, 
---5427, -6380, 4839, 6824, -4212, -7212, 3547, 7538, -2854, -7802, 2134, 7997, -1398, -8127, 648, 8186, 105, -8177, -860, 8097, 1606, -7950, -2340, 7733, 3053, -7452, -3741, 7106, 4397, -6701, 
---5016, 6237, 5591, -5721, -6121, 5155, 6596, -4546, -7017, 3896, 7377, -3215, -7675, 2504, 7906, -1773, -8071, 1026, 8165, -271, -8191, -489, 8145, 1242, -8030, -1987, 7845, 2713, -7595, -3418, 
--7277, 4092, -6899, -4732, 6459, 5331, -5965, -5885, 5418, 6387, -4826, -6836, 4190, 7224, -3520, -7552, 2818, 7813, -2093, -8008, 1348, 8133, -593, -8189, -170, 8172, 929, -8087, -1682, 7929, 
--2419, -7705, -3138, 7412, 3827, -7056, -4485, 6638, 5102, -6163, -5678, 5633, 6202, -5056, -6674, 4433, 7086, -3773, -7439, 3078, 7725, -2358, -7946, 1615, 8096, -860, -8178, 95, 8185, 668, 
---8124, -1428, 7990, 2174, -7787, -2903, 7515, 3605, -7179, -4277, 6778, 4910, -6319, -5503, 5803, 6045, -5238, -6536, 4625, 6968, -3974, -7342, 3285, 7649, -2569, -7890, 1828, 8061, -1074, -8162, 
--307, 8190, 460, -8148, -1226, 8032, 1979, -7847, -2716, 7591, 3428, -7270, -4112, 6883, 4758, -6437, -5364, 5932, 5920, -5376, -6427, 4771, 6874, -4125, -7263, 3441, 7586, -2728, -7844, 1988, 
--8030, -1233, -8147, 465, 8190, 306, -8162, -1076, 8060, 1834, -7888, -2579, 7644, 3299, -7334, -3992, 6956, 4647, -6519, -5263, 6021, 5831, -5471, -6348, 4871, 6807, -4229, -7208, 3547, 7542, 
---2835, -7811, 2096, 8008, -1340, -8136, 569, 8188, 205, -8170, -979, 8076, 1742, -7913, -2492, 7676, 3218, -7372, -3917, 7000, 4580, -6567, -5203, 6073, 5778, -5526, -6302, 4927, 6769, -4286, 
---7176, 3604, 7517, -2892, -7793, 2151, 7996, -1393, -8129, 620, 8187, 157, -8173, -935, 8083, 1702, -7923, -2456, 7688, 3186, -7386, -3890, 7015, 4556, -6582, -5184, 6088, 5762, -5540, -6291, 
--4940, 6760, -4297, -7171, 3613, 7514, -2898, -7791, 2155, 7996, -1393, -8129, 617, 8187, 163, -8173, -944, 8082, 1714, -7919, -2471, 7682, 3204, -7377, -3910, 7003, 4578, -6566, -5206, 6068, 
--5785, -5516, -6313, 4911, 6782, -4263, -7191, 3574, 7532, -2854, -7806, 2106, 8007, -1341, -8136, 560, 8189, 223, -8168, -1007, 8071, 1779, -7901, -2538, 7657, 3271, -7344, -3976, 6962, 4643, 
---6517, -5270, 6011, 5846, -5451, -6370, 4838, 6833, -4183, -7236, 3486, 7570, -2760, -7836, 2006, 8028, -1235, -8148, 450, 8190, 336, -8159, -1122, 8050, 1896, -7868, -2654, 7612, 3386, -7287, 
---4089, 6892, 4752, -6435, -5373, 5916, 5942, -5344, -6459, 4721, 6913, -4055, -7305, 3349, 7627, -2614, -7880, 1853, 8058, -1076, -8163, 287, 8190, 503, -8142, -1291, 8016, 2065, -7818, -2821, 
--7544, 3550, -7202, -4247, 6790, 4903, -6317, -5515, 5782, 6074, -5195, -6578, 4558, 7018, -3879, -7394, 3162, 7700, -2417, -7935, 1647, 8094, -863, -8178, 69, 8184, 723, -8115, -1512, 7967, 
--2284, -7746, -3036, 7451, 3759, -7087, -4448, 6654, 5093, -6160, -5693, 5606, 6236, -5001, -6723, 4346, 7145, -3653, -7501, 2922, 7784, -2166, -7996, 1387, 8130, -596, -8189, -202, 8169, 996, 
---8072, -1784, 7898, 2552, -7650, -3299, 7328, 4012, -6937, -4689, 6479, 5320, -5961, -5903, 5384, 6427, -4758, -6892, 4085, 7290, -3374, -7620, 2629, 7876, -1860, -8059, 1072, 8163, -275, -8191, 
---526, 8138, 1321, -8010, -2105, 7803, 2868, -7523, -3605, 7170, 4306, -6749, -4967, 6262, 5580, -5716, -6140, 5114, 6640, -4464, -7079, 3770, 7447, -3040, -7746, 2280, 7969, -1499, -8117, 702, 
--8185  
--)
--)
-- port map ( 
--			Clk_96 => Clk_96,
--			Ce_F6 => Ce_F6,
--			EN =>EN,
--			Rom_cos_all => Rom_cos_L3_minus--out
--			 );

--P2_PFT <= P2 & PFT;

----  ---
---------------------------------------------------------------------
--MUX_signal_type_cos: process (P2_PFT, Rom_cos_L40_i, Rom_cos_L60_i,
--                                         Rom_cos_L33_i, Rom_cos_L32_i,
--                                         Rom_cos_L22_i, Rom_cos_L21_i, 
--                                        Rom_cos_L16_i, Rom_cos_L15_i,Rom_cos_L23_i )
                                         
--MUX_signal_type_cos: process (PFT,Rom_cos_L23_i ,Rom_cos_L7C3_i)
--
--	begin
--		case PFT is
----		when "0100" => Rom_cos_i <= Rom_cos_L60_i;
----      when "0000" => Rom_cos_i <= Rom_cos_L40_i;
----      when "1001" => Rom_cos_i <= Rom_cos_L33_i;
----		when "0001" => Rom_cos_i <= Rom_cos_L32_i;
----      when "1010" => Rom_cos_i <= Rom_cos_L22_i;
----		when "0010" => Rom_cos_i <= Rom_cos_L21_i;
----      when "1011" => Rom_cos_i <= Rom_cos_L16_i;
----		when "0011" => Rom_cos_i <= Rom_cos_L15_i;
--
--			when "001010" => Rom_cos_i <= Rom_cos_L23_i;
--      --when "001010" => Rom_cos_i <= Rom_cos_L23_i;			
--		
--			when others => Rom_cos_i <= Rom_cos_L23_i;
--      --when others => Rom_cos_i <= Rom_cos_L40_i;
--		              
--		end case;
--end process;

------------------------------------------------------------------------
-------------------------------------------------------------------


----------------------------------------------------------------------
--Converter_cos_sin : process (Clk_96, Ce_F6, NT_PPZ, Sign_LCHM, Rom_cos_i)
--   begin
--       if Clk_96'event and Clk_96 = '1' then
--         if Ce_F6 = '1'  then
--			  if Sign_LCHM = '0'  then
--			      if NT_PPZ = "10001" or NT_PPZ = "10010" or NT_PPZ = "11100" then
--                 -- Rom_cos <= conv_std_logic_vector(-Rom_cos_i, 8);
--                  Rom_cos <= conv_std_logic_vector(-Rom_cos_i, data_rom);
--					else
--						 --Rom_cos <= conv_std_logic_vector(Rom_cos_i, 8);
--						 Rom_cos <= conv_std_logic_vector(Rom_cos_i, data_rom);
--				   end if;
--					
--				elsif Sign_LCHM = '1'  then
--				
--				   if NT_PPZ = "10001" or NT_PPZ = "10010" or NT_PPZ = "11100" then
--                  --Rom_cos <= conv_std_logic_vector(-Rom_cos_i, 8);
--                  Rom_cos <= conv_std_logic_vector(-Rom_cos_i, data_rom);
--                  
--					else 
--						 --Rom_cos <= conv_std_logic_vector(Rom_cos_i, 8);
--						   Rom_cos <= conv_std_logic_vector(Rom_cos_i, data_rom);
--				   end if; 
--				end if;
--			end if; 
--		end if;
--    end process;


	--process (Clk_96, Sign_LCHM, Rom_cos_L3_minus, Rom_cos_L3_plus)
--	begin
--	 if rising_edge(clk_96) then
--    if Sign_LCHM = '1' then
--       Rom_cos_i <= Rom_cos_L3_plus;
--    else
--       Rom_cos_i <= Rom_cos_L3_minus;
--    end if;	
--  end if;	
--   end process;
   
  Rom_cos_i <= Rom_cos_L3_plus when rising_edge(Clk_96);
 ------------------------------------------------------------- 
	process (Clk_96, Ce_F6, EN, Rom_cos_i )
	begin
	  if Clk_96'event and Clk_96 = '1' then
		if Ce_F6 = '1'  then
			if EN = '1' then
				Rom_cos_out <= conv_std_logic_vector(Rom_cos_i, data_rom);
			else
				Rom_cos_out <=(others => '0');
			end if;
		end if;
	  end if;
   end process;

Rom_cos <= Rom_cos_out when rising_edge(Clk_96);

end Behavioral;

