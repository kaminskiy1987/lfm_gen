
--������������� �� ������------ �� �������--------
library IEEE;
	use IEEE.STD_LOGIC_1164.ALL;
	Use ieee.std_logic_arith.all;
	Use ieee.std_logic_unsigned.all;
	USE ieee.math_real.all;
	USE std.textio.ALL;
	USE IEEE.std_logic_textio.ALL;

library elementary;
	use elementary.s274types_pkg.all;
	use elementary.utility.all;
	use elementary.all;
    
entity MUX_signal_type_MP3 is
       generic (
	
	   data_pft: integer := 6;
		data_ppz : integer := 5;
		pft_widht : integer:= 6;
		pft_code : int_array := (10,27);
		data_rom : integer := 12
				);
	Port(
		Clk_96 : in std_logic;
		Ce_F6 : in std_logic;
		En : in std_logic;      
		OD : in std_logic;		
	        LG : in std_logic;		
	        TI : in std_logic;
		PFT : in std_logic_vector (7 downto 0);		
		Sign_LCHM : in std_logic;
		Rom_cos : out std_logic_vector (13 downto 0)		
	);

end MUX_signal_type_MP3;

architecture Behavioral of MUX_signal_type_MP3 is

	signal P2_PFT : std_logic_vector(7 downto 0) := (others => '0');
    signal PFT_adress : std_logic_vector(9 downto 0) := (others => '0');
	signal Rom_cos_i : integer;
	signal adress : std_logic_vector(1 downto 0);  
	signal Rom_cos_L15_i : integer;
	signal Rom_cos_L21_i : integer;
	signal Rom_cos_L32_i : integer;
	signal Rom_cos_L40_i : integer;
begin

    L15_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-7502, 2665, 7936, -1372, -8161, 45, 8167, 1278, -7961, -2566, 7546, 3781, -6939, -4897, 6152, 5883, -5211, -6716, 4138, 7375, -2966, -7847, 1719, 8119, -436, -8189, -857, 8053, 2123, -7720, -3335, 7197, 4460, -6501, -5475, 5648, 6353, -4662, -7077, 3565, 7627, -2389, -7996, 1157, 8173, 96, -8159, -1346, 7953, 2559, -7564, -3710, 7000, 4771, -6278, -5721, 5413, 6537, -4430, -7203, 3348, 7704, -2197, -8034, 997, 8181, 219, -8150, -1428, 7937, 2600, -7555, -3715, 7007, 4743, -6312, -5669, 5483, 6468, -4541, -7130, 3503, 7638, -2398, -7986, 1244, 8164, -69, -8175, -1105, 8016, 2251, -7695, -3349, 7218, 4374, -6598, -5310, 5846, 6135, -4981, -6837, 4019, 7401, -2983, -7819, 1890, 8082, -766, -8189, -371, 8137, 1495, -7931, -2590, 7574, 3630, -7077, -4600, 6447, 5479, -5702, -6255, 4851, 6912, -3917, -7443, 2912, 7834, -1859, -8084, 775, 8187, 317, -8146, -1403, 7959, 2457, -7634, -3467, 7176, 4412, -6597, -5279, 5904, 6050, -5115, -6718, 4240, 7268, -3298, -7696, 2302, 7992, -1274, -8157, 226, 8185, 820, -8081, -1850, 7845, 2846, -7485, -3794, 7005, 4676, -6418, -5483, 5730, 6199, -4956, -6818, 4106, 7328, -3198, -7725, 2243, 8001, -1259, -8156, 257, 8187, 742, -8097, -1729, 7886, 2685, -7562, -3600, 7127, 4457, -6592, -5249, 5963, 5960, -5253, -6587, 4470, 7116, -3628, -7546, 2738, 7867, -1815, -8081, 868, 8181, 84, -8172, -1034, 8052, 1964, -7826, -2867, 7495, 3726, -7070, -4535, 6552, 5279, -5953, -5955, 5278, 6550, -4541, -7062, 3747, 7481, -2912, -7807, 2042, 8033, -1152, -8161, 250, 8188, 649, -8118, -1539, 7949, 2405, -7688, -3241, 7336, 4034, -6901, -4778, 6387, 5462, -5803, -6083, 5154, 6630, -4451, -7103, 3700, 7492, -2913, -7798, 2095, 8017, -1260, -8149, 412, 8190, 434, -8147, -1273, 8015, 2094, -7802, -2891, 7507, 3652, -7138, -4375, 6695, 5048, -6189, -5670, 5621, 6229, -5002, -6727, 4335, 7155, -3630, -7513, 2891, 7795, -2130, -8004, 1351, 8134, -564, -8190, -226, 8167, 1008, -8072, -1780, 7901, 2529, -7663, -3255, 7355, 3946, -6985, -4601, 6554, 5211, -6071, -5775, 5536, 6285, -4958, -6741, 4340, 7137, -3690, -7473, 3012, 7745, -2314, -7954, 1599, 8096, -876, -8175, 149, 8188, 574, -8138, -1291, 8024, 1993, -7851, -2677, 7617, 3336, -7330, -3968, 6988, 4566, -6599, -5130, 6162, 5652, -5685, -6132, 5168, 6565, -4620, -6951, 4041, 7286, -3439, -7570, 2815, 7800, -2177, -7979, 1527, 8102, -872, -8174, 213, 8190, 441, -8155, -1091, 8068, 1729, -7933, -2354, 7747, 2959, -7517, -3544, 7242, 4103, -6926, -4636, 6570, 5137, -6180, -5608, 5754, 6041, -5301, -6440, 4818, 6798, -4313, -7119, 3786, 7397, -3244, -7636, 2686, 7830, -2119, -7984, 1542, 8094, -963, -8164, 381, 8190, 197, -8177, -773, 8122, 1339, -8030, -1897, 7898, 2440, -7731, -2970, 7528, 3481, -7293, -3975, 7024, 4445, -6728, -4894, 6402, 5317, -6052, -5716, 5677, 6086, -5282, -6429, 4866, 6741, -4434, -7026, 3986, 7278, -3526, -7501, 3055, 7691, -2576, -7852, 2089, 7980, -1600, -8079, 1107, 8145, -615, -8183, 122, 8190, 365, -8169, -849, 8118, 1324, -8042, -1794, 7937, 2251, -7808, -2700, 7653, 3134, -7476, -3557, 7275, 3964, -7055, -4356, 6814, 4730, -6555, -5089, 6277, 5428, -5986, -5751, 5677, 6052, -5357, -6336, 5023, 6598, -4680, -6842, 4326, 7063, -3965, -7267, 3596, 7447, -3222, -7610, 2842, 7750, -2460, -7872, 2074, 7972, -1688, -8054, 1300, 8115, -915, -8160, 530, 8183, -149, -8191, -230, 8180, 604, -8153, -974, 8108, 1337, -8050, -1695, 7974, 2045, -7886, -2388, 7781, 2722, -7666, -3050, 7536, 3366, -7396, -3675, 7242, 3973, -7081, -4262, 6907, 4540, -6726, -4809, 6534, 5065, -6337, -5313, 6130, 5548, -5919, -5774, 5700, 5988, -5477, -6192, 5247, 6383, -5016, -6566, 4779, 6736, -4540, -6897, 4297, 7046, -4054, -7187, 3808, 7315, -3562, -7435, 3314, 7544, -3067, -7645, 2819, 7734, -2573, -7817, 2326, 7888, -2082, -7953, 1839, 8008, -1599, -8057, 1359, 8096, -1124, -8129, 889, 8154, -660, -8173, 431, 8184, -208, -8191, -13, 8190, 229, -8185, -443, 8172, 650, -8157, -856, 8134, 1056, -8110, -1253, 8079, 1443, -8046, -1632, 8007, 1814, -7967, -1993, 7922, 2165, -7876, -2335, 7826, 2499, -7775, -2660, 7720, 2814, -7665, -2965, 7606, 3110, -7548, -3253, 7487, 3389, -7427, -3522, 7364, 3649, -7302, -3773, 7238, 3892, -7176, -4007, 7112, 4117, -7050, -4225, 6986, 4326, -6925, -4425, 6862, 4518, -6802, -4610, 6741, 4695, -6682, -4779, 6623, 4857, -6567, -4933, 6511, 5004, -6458, -5073, 6405, 5137, -6355, -5199, 6305, 5256, -6259, -5312, 6213, 5363, -6170, -5412, 6128, 5456, -6090, -5499, 6052, 5537, -6019, -5575, 5985, 5607, -5956, -5638, 5928, 5665, -5904, -5691, 5880, 5712, -5861, -5732, 5843, 5748, -5829, -5763, 5815, 5773, -5806, -5782, 5798, 5787, -5794, -5792, 5791, 5791, -5793, -5790, 5795, 5785, -5802, -5779, 5810, 5768, -5822, -5756, 5835, 5740, -5852, -5723, 5870, 5701, -5892, -5679, 5915, 5652, -5942, -5624, 5970, 5591, -6002, -5557, 6035, 5518, -6071, -5479, 6108, 5434, -6149, -5388, 6191, 5337, -6236, -5285, 6281, 5228, -6330, -5169, 6379, 5105, -6432, -5040, 6484, 4969, -6540, -4896, 6595, 4818, -6653, -4738, 6711, 4653, -6772, -4565, 6831, 4472, -6894, -4377, 6955, 4275, -7018, -4172, 7080, 4062, -7144, -3951, 7207, 3833, -7271, -3712, 7333, 3585, -7396, -3456, 7457, 3321, -7518, -3182, 7577, 3038, -7636, -2891, 7692, 2737, -7748, -2580, 7800, 2417, -7852, -2251, 7899, 2079, -7946, -1904, 7987, 1723, -8027, -1539, 8062, 1348, -8095, -1155, 8122, 956, -8147, -754, 8165, 547, -8180, -337, 8187, 121, -8191, 97, 8188, -320, -8180, 544, 8164, -774, -8143, 1005, 8113, -1241, -8078, 1478, 8033, -1719, -7982, 1960, 7921, -2205, -7854, 2449, 7776, -2696, -7691, 2942, 7595, -3191, -7491, 3437, 7376, -3685, -7252, 3931, 7117, -4176, -6973, 4418, 6817, -4660, -6653, 4897, 6476, -5133, -6289, 5362, 6091, -5589, -5883, 5809, 5662, -6026, -5433, 6234, 5190, -6437, -4939, 6631, 4675, -6818, -4403, 6994, 4118, -7163, -3826, 7320, 3521, -7468, -3210, 7602, 2887, -7726, -2557, 7835, 2217, -7932, -1871, 8013, 1516, -8082, -1157, 8132, 789, -8169, -418, 8187, 41, -8190, 339, 8173, -723, -8140, 1107, 8087, -1495, -8016, 1881, 7924, -2268, -7814, 2651, 7682, -3033, -7531, 3409, 7359, -3782, -7168, 4146, 6955, -4505, -6723, 4853, 6469, -5192, -6197, 5518, 5903, -5834, -5593, 6133, 5261, -6419, -4913, 6686, 4545, -6937, -4162, 7167, 3762, -7379, -3348, 7567, 2918, -7734, -2478, 7875, 2023, -7993, -1561, 8083, 1087, -8147, -608, 8182, 121, -8191, 368, 8167, -861, -8116, 1353, 8033, -1846, -7920, 2333, 7775, -2817, -7600, 3291, 7393, -3758, -7156, 4211, 6887, -4652, -6589, 5075, 6260, -5482, -5905, 5867, 5519, -6231, -5110, 6568, 4672, -6880, -4213, 7162, 3730, -7415, -3229, 7633, 2707, -7819, -2171, 7968, 1619, -8081, -1057, 8154, 485, -8189, 91, 8182, -673, -8135, 1253, 8044, -1832, -7913, 2403, 7738, -2967, -7522, 3517, 7263, -4053, -6964, 4568, 6623, -5063, -6246, 5531, 5828, -5972, -5377, 6379, 4890, -6753, -4374, 7089, 3826, -7385, -3255, 7637, 2658, -7846, -2044, 8006, 1411, -8119, -768, 8179, 114, -8189, 542, 8144, -1201, -8048, 1853, 7896, -2498, -7692, 3128, 7434, -3743, -7125, 4333, 6764, -4899, -6355, 5431, 5897, -5929, -5396, 6385, 4853, -6800, -4272, 7165, 3656, -7481, -3010, 7741, 2337, -7945, -1645, 8088, 934, -8171, -214, 8189, -513, -8145, 1238, 8033, -1958, -7858, 2664, 7617, -3354, -7313, 4018, 6946, -4654, -6521, 5252, 6036, -5810, -5500, 6319, 4911, -6777, -4279, 7177, 3604, -7517, -2896, 7790, 2157, -7996, -1396, 8128, 618, -8188, 169, 8171, -959, -8079, 1742, 7909, -2514, -7664, 3264, 7343, -3987, -6950, 4673, 6486, -5318, -5958, 5912, 5365, -6451, -4719, 6924, 4019, -7332, -3277, 7664, 2495, -7919, -1687, 8091, 854, -8180, -12, 8180, -837, -8094, 1679, 7918, -2507, -7656, 3310, 7307, -4081, -6877, 4809, 6365, -5486, -5782, 6103, 5127, -6654, -4413, 7128, 3643, -7523, -2828, 7829, 1975, -8046, -1097, 8165, 200, -8188, 701, 8109, -1600, -7933, 2480, 7656, -3335, -7284, 4150, 6817, -4918, -6264, 5624, 5626, -6263, -4916, 6821, 4137, -7295, -3302, 7673, 2419, -7952, -1502, 8125, 560, -8191, 392, 8144, -1344, -7988, 2279, 7719, -3189, -7344, 4055, 6863, -4870, -6286, 5617, 5614, -6289, -4863, 6871, 4036, -7358, -3149, 7738, 2211, -8007, -1239, 8157, 243, -8187, 759, 8093, -1754, -7878, 2725, 7540, -3660, -7088, 4539, 6521, -5353, -5854, 6085, 5089, -6725, -4244, 7259, 3326, -7681, -2354, 7979, 1338, -8150, -298, 8187, -752, -8092, 1791, 7860, -2806, -7498, 3776, 7008, -4687, -6399, 5520, 5677, -6264, -4857, 6901, 3948, -7422, -2970, 7813, 1934, -8071, -863, 8184, -229, -8155, 1319, 7977, -2391, -7656, 3421, 7194, -4394, -6600, 5288, 5881, -6089, -5052, 6777, 4124, -7343, -3118, 7770, 2047, -8054, -936, 8182, -198, -8156, 1331, 7969, -2443, -7629, 3509, 7136, -4512, -6503, 5426, 5737, -6237, -4855, 6924, 3871, -7476, -2808, 7875, 1682, -8117, -520, 8190, -658, -8096, 1825, 7832, -2959, -7404, 4032, 6817, -5025, -6086, 5913, 5220, -6678, -4241, 7300, 3166, -7768, -2021, 8065, 826, -8189, 389, 8130, -1601, -7892, 2779, 7475, -3900, -6890, 4935, 6146, -5863, -5262, 6657, 4253, -7303, -3144, 7780, 1958, -8080, -724, 8190, -532, -8109, 1777, 7835, -2986, -7375, 4125, 6735, -5171, -5933, 6092, 4983, -6870, -3911, 7481, 2738, -7911, -1496, 8146, 211, -8180, 1080, 8008, -2350, -7636, 3562, 7068, -4690, -6320, 5699, 5407, -6566, -4354, 7265, 3184, -7779, -1929, 8090, 619, -8191, 710, 8075, -2025, -7746) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L15_i
    );

    L21_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-5863, 5222, 6715, -4127, -7388, 2924, 7863, -1647, -8131, 327, 8184, 997, -8023, -2294, 7652, 3527, -7085, -4668, 6334, 5684, -5423, -6554, 4372, 7253, -3214, -7767, 1974, 8081, -689, -8191, -614, 8093, 1896, -7794, -3130, 7298, 4282, -6623, -5327, 5784, 6236, -4805, -6991, 3707, 7571, -2523, -7967, 1278, 8165, -6, -8167, -1266, 7970, 2502, -7582, -3678, 7012, 4761, -6278, -5731, 5393, 6561, -4385, -7235, 3273, 7737, -2089, -8057, 856, 8187, 392, -8128, -1631, 7879, 2827, -7451, -3958, 6851, 4994, -6097, -5916, 5204, 6699, -4196, -7331, 3094, 7794, -1926, -8084, 716, 8190, 505, -8115, -1715, 7859, 2883, -7432, -3986, 6841, 4998, -6103, -5900, 5231, 6670, -4250, -7296, 3177, 7762, -2041, -8061, 860, 8186, 334, -8139, -1520, 7917, 2670, -7530, -3763, 6984, 4773, -6295, -5682, 5474, 6470, -4544, -7125, 3520, 7629, -2428, -7977, 1286, 8160, -123, -8179, -1042, 8029, 2182, -7721, -3277, 7256, 4302, -6650, -5241, 5910, 6072, -5057, -6783, 4104, 7358, -3075, -7789, 1987, 8065, -864, -8186, -276, 8147, 1405, -7953, -2507, 7606, 3556, -7116, -4538, 6491, 5429, -5746, -6218, 4894, 6887, -3953, -7428, 2940, 7827, -1876, -8083, 778, 8187, 330, -8144, -1431, 7950, 2502, -7614, -3527, 7139, 4484, -6539, -5360, 5822, 6136, -5004, -6804, 4098, 7348, -3124, -7763, 2095, 8039, -1034, -8177, -45, 8170, 1118, -8024, -2172, 7738, 3183, -7323, -4140, 6783, 5023, -6130, -5820, 5374, 6516, -4532, -7102, 3614, 7568, -2640, -7908, 1623, 8116, -584, -8191, -465, 8131, 1501, -7941, -2512, 7621, 3478, -7181, -4388, 6625, 5224, -5967, -5977, 5214, 6631, -4383, -7181, 3483, 7616, -2533, -7933, 1544, 8124, -536, -8191, -480, 8131, 1484, -7949, -2465, 7644, 3404, -7227, -4292, 6701, 5111, -6077, -5853, 5363, 6505, -4573, -7061, 3716, 7510, -2809, -7851, 1861, 8074, -891, -8182, -92, 8170, 1069, -8043, -2030, 7800, 2957, -7450, -3843, 6993, 4670, -6442, -5431, 5801, 6114, -5082, -6712, 4294, 7214, -3451, -7618, 2561, 7915, -1641, -8107, 700, 8187, 247, -8160, -1190, 8022, 2112, -7780, -3006, 7435, 3856, -6995, -4655, 6463, 5390, -5851, -6055, 5164, 6639, -4414, -7138, 3609, 7544, -2762, -7855, 1880, 8064, -980, -8175, 67, 8181, 841, -8089, -1739, 7896, 2610, -7608, -3450, 7228, 4243, -6763, -4985, 6217, 5664, -5600, -6275, 4916, 6808, -4179, -7261, 3392, 7627, -2571, -7905, 1720, 8089, -854, -8181, -22, 8178, 893, -8084, -1753, 7897, 2588, -7624, -3395, 7265, 4159, -6829, -4877, 6316, 5537, -5738, -6137, 5098, 6667, -4406, -7125, 3667, 7503, -2893, -7803, 2089, 8016, -1267, -8147, 432, 8190, 402, -8150, -1232, 8024, 2045, -7818, -2836, 7531, 3594, -7171, -4315, 6737, 4989, -6240, -5612, 5679, 6176, -5067, -6680, 4404, 7114, -3703, -7480, 2966, 7771, -2205, -7988, 1423, 8126, -633, -8188, -164, 8171, 954, -8080, -1735, 7912, 2495, -7674, -3231, 7363, 3934, -6989, -4600, 6551, 5221, -6057, -5795, 5509, 6314, -4915, -6777, 4279, 7176, -3609, -7514, 2908, 7784, -2186, -7987, 1445, 8120, -697, -8185, -56, 8179, 804, -8107, -1545, 7965, 2269, -7760, -2973, 7490, 3649, -7162, -4295, 6775, 4902, -6337, -5469, 5848, 5989, -5316, -6462, 4743, 6881, -4136, -7246, 3498, 7552, -2836, -7802, 2154, 7988, -1460, -8116, 755, 8181, -49, -8186, -657, 8128, 1353, -8014, -2039, 7839, 2705, -7610, -3352, 7325, 3970, -6991, -4559, 6607, 5113, -6180, -5630, 5710, 6104, -5203, -6537, 4661, 6921, -4092, -7259, 3494, 7544, -2878, -7780, 2243, 7962, -1597, -8092, 942, 8167, -285, -8191, -373, 8161, 1025, -8080, -1669, 7946, 2298, -7765, -2913, 7535, 3505, -7261, -4074, 6941, 4615, -6583, -5128, 6184, 5606, -5752, -6050, 5285, 6455, -4792, -6822, 4270, 7146, -3728, -7430, 3165, 7668, -2588, -7864, 1997, 8012, -1399, -8118, 794, 8176, -189, -8191, -416, 8159, 1015, -8086, -1607, 7967, 2187, -7810, -2754, 7609, 3302, -7372, -3833, 7096, 4340, -6787, -4825, 6443, 5281, -6071, -5711, 5667, 6108, -5240, -6476, 4786, 6809, -4314, -7109, 3821, 7372, -3314, -7601, 2792, 7791, -2261, -7946, 1720, 8061, -1176, -8142, 627, 8183, -80, -8189, -467, 8157, 1008, -8091, -1543, 7989, 2067, -7854, -2582, 7685, 3082, -7486, -3568, 7254, 4034, -6996, -4484, 6708, 4911, -6396, -5319, 6058, 5701, -5699, -6060, 5318, 6392, -4920, -6699, 4503, 6977, -4073, -7229, 3627, 7451, -3173, -7645, 2707, 7809, -2235, -7945, 1756, 8049, -1274, -8126, 789, 8172, -306, -8191, -178, 8180, 657, -8142, -1133, 8076, 1600, -7984, -2062, 7864, 2512, -7722, -2953, 7553, 3381, -7362, -3798, 7148, 4198, -6914, -4584, 6658, 4953, -6385, -5306, 6092, 5639, -5785, -5956, 5460, 6251, -5123, -6528, 4771, 6783, -4410, -7018, 4036, 7231, -3655, -7425, 3264, 7594, -2869, -7745, 2467, 7871, -2062, -7978, 1652, 8062, -1243, -8126, 831, 8167, -421, -8189, 11, 8188, 394, -8170, -798, 8130, 1196, -8072, -1590, 7994, 1976, -7900, -2356, 7786, 2727, -7657, -3091, 7510, 3444, -7349, -3789, 7172, 4121, -6982, -4445, 6776, 4755, -6560, -5054, 6329, 5340, -6090, -5614, 5838, 5873, -5578, -6121, 5307, 6354, -5029, -6574, 4742, 6779, -4451, -6971, 4151, 7147, -3848, -7311, 3538, 7459, -3227, -7595, 2910, 7715, -2592, -7822, 2271, 7914, -1950, -7994, 1627, 8058, -1305, -8111, 982, 8149, -662, -8176, 342, 8188, -26, -8190, -290, 8178, 601, -8157, -910, 8121, 1214, -8077, -1515, 8020, 1810, -7955, -2101, 7877, 2386, -7792, -2666, 7696, 2939, -7593, -3208, 7479, 3469, -7359, -3725, 7230, 3972, -7095, -4214, 6951, 4448, -6803, -4676, 6647, 4895, -6487, -5108, 6319, 5312, -6149, -5511, 5972, 5700, -5792, -5883, 5607, 6057, -5420, -6225, 5228, 6384, -5035, -6537, 4837, 6681, -4639, -6819, 4438, 6948, -4236, -7072, 4032, 7186, -3828, -7296, 3621, 7396, -3416, -7492, 3209, 7579, -3004, -7661, 2796, 7735, -2592, -7804, 2385, 7866, -2182, -7923, 1978, 7972, -1777, -8018, 1575, 8056, -1377, -8091, 1179, 8119, -985, -8143, 790, 8161, -600, -8176, 410, 8184, -224, -8190, 39, 8190, 142, -8188, -322, 8180, 497, -8171, -672, 8155, 841, -8139, -1010, 8117, 1174, -8095, -1336, 8067, 1494, -8039, -1650, 8007, 1802, -7974, -1952, 7936, 2097, -7899, -2240, 7858, 2379, -7817, -2516, 7773, 2648, -7729, -2779, 7681, 2905, -7635, -3030, 7585, 3149, -7537, -3267, 7486, 3380, -7436, -3492, 7383, 3599, -7332, -3705, 7279, 3805, -7227, -3905, 7174, 4000, -7122, -4094, 7068, 4182, -7017, -4270, 6963, 4353, -6913, -4436, 6860, 4513, -6810, -4590, 6759, 4662, -6710, -4734, 6660, 4800, -6613, -4867, 6565, 4928, -6520, -4990, 6473, 5046, -6430, -5103, 6386, 5155, -6345, -5206, 6303, 5253, -6265, -5300, 6226, 5343, -6190, -5386, 6154, 5424, -6121, -5462, 6088, 5496, -6058, -5530, 6028, 5560, -6001, -5590, 5974, 5616, -5951, -5642, 5927, 5664, -5907, -5686, 5887, 5704, -5870, -5722, 5853, 5736, -5840, -5751, 5827, 5761, -5818, -5772, 5808, 5779, -5802, -5785, 5796, 5789, -5794, -5792, 5791, 5791, -5793, -5791, 5794, 5787, -5799, -5783, 5804, 5775, -5813, -5767, 5822, 5756, -5834, -5744, 5846, 5729, -5862, -5714, 5878, 5695, -5897, -5676, 5916, 5653, -5939, -5630, 5962, 5603, -5988, -5576, 6014, 5545, -6043, -5514, 6072, 5479, -6105, -5444, 6137, 5405, -6172, -5365, 6207, 5322, -6246, -5278, 6284, 5230, -6325, -5181, 6365, 5128, -6408, -5075, 6451, 5018, -6497, -4960, 6542, 4897, -6589, -4834, 6636, 4767, -6686, -4699, 6734, 4626, -6785, -4553, 6835, 4474, -6887, -4395, 6937, 4312, -6991, -4227, 7042, 4138, -7096, -4048, 7147, 3952, -7201, -3856, 7253, 3755, -7306, -3653, 7357, 3545, -7410, -3437, 7460, 3324, -7512, -3209, 7561, 3089, -7611, -2968, 7658, 2842, -7706, -2715, 7750, 2582, -7796, -2449, 7837, 2310, -7879, -2169, 7917, 2024, -7956, -1878, 7990, 1726, -8024, -1573, 8053, 1415, -8082, -1256, 8106, 1092, -8129, -926, 8147, 756, -8164, -585, 8175, 409, -8185, -233, 8189, 51, -8191, 131, 8187, -317, -8181, 504, 8169, -695, -8153, 887, 8131, -1082, -8106, 1277, 8074, -1477, -8038, 1675, 7996, -1878, -7949, 2079, 7895, -2284, -7836, 2488, 7770, -2694, -7699, 2899, 7620, -3107, -7537, 3312, 7444, -3519, -7347, 3724, 7241, -3930, -7130, 4134, 7010, -4338, -6885, 4538, 6750, -4739, -6610, 4936, 6461, -5132, -6306, 5324, 6141, -5514, -5971, 5699, 5792, -5883, -5607, 6060, 5412, -6235, -5212, 6403, 5002, -6568, -4787, 6725, 4562, -6878, -4332, 7023, 4094, -7164, -3850, 7295, 3597, -7420, -3340, 7536, 3074, -7646, -2804, 7744, 2526, -7836, -2245, 7917, 1956, -7989, -1663, 8049, 1364, -8101, -1063, 8140, 756, -8169, -446, 8185, 132, -8191, 183, 8183, -502, -8165, 822, 8131, -1144, -8087, 1466, 8027, -1789, -7956, 2110, 7869, -2432, -7771, 2751, 7656, -3069, -7529, 3382, 7387, -3694, -7232, 4000, 7060, -4302, -6877, 4597, 6678, -4887, -6466, 5168, 6239, -5444, -5999, 5708, 5745, -5966, -5479, 6211, 5198, -6447, -4906, 6669, 4601, -6881, -4285, 7078, 3956, -7263, -3618, 7431, 3268, -7586, -2911, 7723, 2542, -7845, -2167, 7949, 1783, -8036, -1394, 8103, 997, -8153, -597, 8181, 191, -8191, 215, 8180, -626, -8149, 1036, 8096, -1448, -8023, 1857, 7927, -2265, -7811, 2668, 7672, -3068, -7513, 3460, 7330, -3847, -7128, 4223, 6903, -4592, -6658, 4948, 6391, -5293, -6106, 5623, 5799, -5941, -5475, 6240, 5131, -6524, -4771, 6788, 4392, -7034, -4000, 7257, 3591, -7461, -3169, 7640, 2734, -7797, -2289, 7927, 1831, -8034, -1368, 8112, 895, -8165, -418, 8189, -64, -8186, 547, 8152, -1032, -8092, 1515, 8000, -1996, -7881, 2471, 7730, -2941, -7552, 3401, 7343, -3852, -7107, 4289, 6841, -4714, -6550, 5121, 6229, -5512, -5884, 5881, 5512, -6230, -5118, 6554, 4700, -6855, -4262, 7128, 3803, -7374, -3327, 7589, 2833, -7774, -2327, 7925, 1806, -8045, -1277, 8128, 738, -8178, -195, 8190, -354, -8167, 901, 8106, -1449, -8009, 1991, 7872, -2528, -7701, 3054, 7490, -3570, -7245, 4069, 6963, -4553, -6647, 5015, 6296, -5457, -5914, 5872, 5499, -6261, -5057, 6619, 4585, -6947, -4090, 7238, 3570, -7496, -3031, 7714, 2472, -7894, -1899, 8031, 1312, -8128, -717, 8180, 113, -8189, 491, 8152, -1097, -8071, 1698, 7943, -2294, -7772, 2878, 7554, -3449, -7294, 4001, 6989, -4534, -6644, 5041, 6257, -5523, -5833, 5972, 5370, -6388, -4876, 6766, 4348, -7107, -3793, 7403, 3211, -7656, -2608, 7861, 1985, -8020, -1349, 8126, 700, -8183, -45, 8186, -614, -8137, 1270, 8033, -1922, -7878, 2562, 7668, -3189, -7408, 3796, 7096, -4381, -6735, 4936, 6326, -5462, -5873, 5949, 5376, -6400, -4841, 6805, 4268, -7165, -3665, 7474, 3031, -7732, -2375, 7933, 1697, -8079, -1006, 8164, 304, -8191, 402, 8156, -1109, -8060, 1808, 7902, -2498, -7685, 3169, 7406, -3821, -7071, 4443, 6678, -5034, -6232, 5587, 5735, -6099, -5191, 6562, 4603, -6976, -3977, 7333, 3314, -7633, -2625, 7870, 1909, -8045, -1177, 8151, 430, -8191, 320, 8161, -1073, -8063, 1817, 7894, -2550, -7658, 3261, 7353, -3948, -6985, 4601, 6552, -5218, -6062, 5789, 5514, -6311, -4917, 6777, 4272, -7185, -3587, 7526, 2866, -7802, -2118, 8005, 1346, -8136, -560, 8189, -235, -8167, 1028, 8066, -1817, -7889, 2588, 7634, -3339, -7307, 4058, 6905, -4742, -6437, 5379, 5901, -5967, -5308, 6496, 4657, -6963, -3960, 7360, 3219, -7685, -2444, 7931, 1640, -8098, -819, 8181, -15, -8180, 850, 8092, -1680, -7921, 2493, 7663, -3285, -7325, 4041, 6905, -4759, -6411, 5425, 5845, -6036, -5215, 6581, 4524, -7057, -3783, 7454, 2995, -7772, -2174, 8001, 1324, -8143, -459, 8190, -417, -8147, 1288, 8008, -2149, -7778, 2985, 7455, -3791, -7046, 4553, 6551, -5266, -5979, 5916, 5332, -6500, -4622, 7005, 3852, -7430, -3035, 7763, 2178, -8005, -1293, 8147, 387, -8191, 524, 8132, -1432, -7973, 2324, 7711, -3190, -7353, 4017, 6899, -4797, -6358, 5516, 5732, -6168, -5032, 6739, 4262, -7227, -3437, 7619, 2563, -7914, -1654, 8104, 719, -8188, 226, 8161, -1173, -8025, 2104, 7780, -3012, -7429, 3879, 6974, -4697, -6424, 5450, 5782, -6132, -5060, 6729, 4263, -7235, -3407, 7638, 2498, -7936, -1553, 8120, 581, -8191, 399, 8142, -1378, -7977, 2338, 7694, -3269, -7300, 4151, 6795, -4977, -6191, 5730, 5492, -6401, -4711, 6976, 3855, -7450, -2941, 7811, 1978, -8056, -985, 8176, -28, -8174, 1041, 8044, -2043, -7790, 3013, 7413, -3941, -6920, 4807, 6316, -5602, -5612, 6308, 4815, -6917, -3942, 7415, 3001, -7797, -2011, 8052, 984, -8178, 59, 8170, -1106, -8029, 2135, 7754, -3134, -7351, 4081, 6823, -4964, -6181, 5764, 5433, -6470, -4592, 7067, 3669, -7547, -2684, 7897, 1648, -8115, -584, 8190, -496, -8126, 1567, 7918, -2615, -7573, 3618, 7091, -4562, -6485, 5424, 5761, -6195, -4934, 6854, 4014, -7394, -3022, 7799, 1971, -8066, -884, 8184, -224, -8154, 1329, 7973, -2413, -7646, 3454, 7174, -4434, -6569, 5332, 5837, -6133, -4996, 6819, 4056, -7379, -3039, 7798, 1960, -8070, -843, 8186, -295, -8146, 1428, 7946, -2537, -7592, 3598, 7088, -4592, -6444, 5496, 5670, -6296, -4784, 6970, 3799, -7508, -2737, 7895, 1616, -8125, -461, 8190, -707, -8090, 1861, 7823, -2982, -7396, 4042, 6815, -5023, -6093, 5899, 5241, -6657, -4280, 7275, 3225, -7744, -2101, 8048, 929, -8185, 263, 8145, -1455, -7933, 2615, 7549, -3724, -7003, 4753, 6302, -5683, -5464, 6489, 4504, -7157, -3445, 7666, 2305, -8010, -1114, 8175, -106, -8160, 1324, 7961, -2517, -7584, 3655, 7034, -4713, -6326, 5666, 5470, -6493, -4490, 7171, 3402, -7688, -2236, 8027, 1014, -8182, 232, 8146, -1477, -7921, 2688, 7508, -3841, -6919, 4903, 6164, -5853, -5262, 6664, 4232, -7320, -3100, 7799, 1889, -8093, -632, 8190, -644, -8091, 1906, 7792, -3125, -7304, 4268, 6634, -5311, -5800, 6222, 4819, -6983, -3719, 7569, 2521, -7969, -1260, 8168, -38, -8163, 1335, 7949, -2603, -7535, 3805, 6926, -4914, -6140, 5897, 5193, -6732, -4111, 7392, 2920, -7864, -1651, 8130, 336, -8185, 989, 8023, -2293, -7652, 3537, 7075, -4691, -6311) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L21_i
    );

    L32_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-8041, -2217, 7678, 3470, -7113, -4630, 6357, 5664, -5437, -6549, 4372, 7258, -3195, -7777, 1933, 8089, -625, -8191, -700, 8077, 2003, -7755, -3255, 7230, 4418, -6520, -5467, 5640, 6372, -4618, -7114, 3477, 7670, -2250, -8031, 966, 8184, 340, -8131, -1638, 7869, 2890, -7410, -4069, 6763, 5142, -5948, -6087, 4982, 6875, -3895, -7492, 2710, 7919, -1460, -8150, 175, 8177, 1112, -8003, -2371, 7630, 3568, -7071, -4678, 6337, 5669, -5450, -6523, 4430, 7214, -3305, -7730, 2099, 8056, -846, -8189, -428, 8121, 1688, -7861, -2907, 7409, 4053, -6783, -5103, 5994, 6028, -5065, -6809, 4015, 7427, -2873, -7869, 1663, 8124, -417, -8189, -839, 8059, 2071, -7744, -3255, 7246, 4360, -6582, -5364, 5764, 6240, -4816, -6973, 3756, 7542, -2613, -7939, 1410, 8152, -178, -8180, -1059, 8019, 2267, -7678, -3424, 7162, 4501, -6486, -5476, 5664, 6324, -4717, -7032, 3664, 7579, -2532, -7958, 1343, 8157, -129, -8177, -1089, 8014, 2279, -7677, -3419, 7169, 4481, -6506, -5445, 5700, 6286, -4773, -6991, 3741, 7542, -2632, -7930, 1465, 8144, -270, -8185, -931, 8048, 2108, -7740, -3240, 7266, 4300, -6640, -5269, 5871, 6123, -4982, -6848, 3986, 7425, -2910, -7848, 1773, 8104, -602, -8191, -582, 8107, 1750, -7855, -2882, 7440, 3950, -6873, -4938, 6164, 5821, -5331, -6585, 4389, 7211, -3360, -7692, 2262, 8013, -1122, -8174, -41, 8167, 1200, -7998, -2335, 7666, 3419, -7183, -4435, 6556, 5360, -5801, -6178, 4930, 6871, -3965, -7429, 2921, 7838, -1823, -8094, 689, 8190, 454, -8127, -1590, 7905, 2690, -7531, -3739, 7010, 4712, -6357, -5595, 5581, 6367, -4701, -7018, 3730, 7532, -2692, -7904, 1602, 8123, -485, -8191, -641, 8102, 1751, -7863, -2828, 7475, 3849, -6951, -4799, 6295, 5656, -5526, -6409, 4653, 7040, -3698, -7543, 2675, 7905, -1606, -8123, 507, 8190, 597, -8111, -1690, 7882, 2750, -7514, -3760, 7009, 4698, -6380, -5553, 5636, 6306, -4795, -6947, 3868, 7461, -2875, -7845, 1832, 8087, -760, -8189, -326, 8145, 1403, -7960, -2455, 7635, 3461, -7180, -4407, 6599, 5274, -5908, -6050, 5113, 6719, -4234, -7274, 3283, 7702, -2279, -8000, 1235, 8160, -175, -8184, -889, 8067, 1934, -7818, -2947, 7436, 3907, -6932, -4802, 6312, 5615, -5590, -6334, 4776, 6947, -3885, -7446, 2931, 7820, -1932, -8068, 901, 8182, 141, -8165, -1181, 8014, 2198, -7736, -3180, 7332, 4107, -6813, -4969, 6185, 5749, -5461, -6437, 4650, 7021, -3769, -7495, 2827, 7849, -1845, -8081, 834, 8184, 186, -8162, -1204, 8011, 2200, -7738, -3162, 7345, 4071, -6842, -4919, 6233, 5688, -5531, -6372, 4745, 6955, -3891, -7434, 2977, 7798, -2022, -8047, 1036, 8173, -38, -8178, -960, 8061, 1941, -7825, -2893, 7473, 3799, -7014, -4649, 6450, 5428, -5795, -6129, 5055, 6737, -4245, -7248, 3373, 7653, -2456, -7948, 1503, 8127, -532, -8191, -446, 8137, 1414, -7970, -2363, 7688, 3275, -7301, -4141, 6810, 4945, -6226, -5682, 5555, 6335, -4810, -6902, 3998, 7371, -3134, -7739, 2226, 7999, -1292, -8151, 340, 8189, 613, -8119, -1558, 7937, 2478, -7651, -3366, 7260, 4204, -6775, -4987, 6199, 5701, -5544, -6339, 4814, 6891, -4025, -7353, 3182, 7717, -2301, -7980, 1390, 8138, -464, -8191, -467, 8138, 1390, -7981, -2294, 7721, 3166, -7364, -3997, 6913, 4775, -6376, -5492, 5759, 6138, -5072, -6706, 4321, 7188, -3519, -7582, 2674, 7879, -1798, -8079, 900, 8178, 5, -8179, -910, 8077, 1801, -7880, -2670, 7585, 3503, -7201, -4294, 6729, 5030, -6180, -5707, 5555, 6312, -4868, -6843, 4123, 7291, -3332, -7653, 2502, 7923, -1645, -8102, 770, 8184, 111, -8173, -991, 8066, 1855, -7868, -2699, 7578, 3508, -7204, -4278, 6747, 4995, -6217, -5657, 5615, 6252, -4954, -6777, 4236, 7224, -3475, -7591, 2674, 7871, -1848, -8066, 1001, 8170, -146, -8187, -710, 8112, 1555, -7951, -2383, 7702, 3182, -7373, -3947, 6963, 4666, -6482, -5336, 5931, 5946, -5320, -6494, 4652, 6970, -3939, -7375, 3184, 7699, -2399, -7944, 1589, 8105, -766, -8184, -65, 8176, 891, -8087, -1709, 7914, 2506, -7663, -3278, 7332, 4013, -6931, -4708, 6459, 5352, -5926, -5944, 5332, 6474, -4690, -6941, 4000, 7336, -3275, -7661, 2517, 7909, -1738, -8081, 943, 8173, -141, -8187, -662, 8122, 1454, -7981, -2234, 7762, 2988, -7473, -3715, 7111, 4403, -6686, -5050, 6198, 5647, -5654, -6192, 5058, 6677, -4418, -7102, 3738, 7458, -3026, -7748, 2287, 7965, -1530, -8111, 760, 8182, 14, -8182, -788, 8106, 1551, -7961, -2301, 7744, 3026, -7462, -3726, 7112, 4389, -6704, -5015, 6236, 5594, -5717, -6125, 5149, 6601, -4539, -7021, 3890, 7379, -3212, -7675, 2506, 7904, -1783, -8068, 1045, 8163, -301, -8191, -445, 8150, 1184, -8043, -1913, 7869, 2623, -7634, -3312, 7334, 3971, -6979, -4598, 6566, 5185, -6103, -5731, 5591, 6228, -5038, -6677, 4444, 7070, -3819, -7409, 3163, 7687, -2487, -7907, 1791, 8063, -1084, -8159, 369, 8190, 345, -8161, -1057, 8069, 1757, -7917, -2444, 7705, 3109, -7437, -3751, 7113, 4362, -6739, -4942, 6315, 5481, -5847, -5982, 5336, 6435, -4789, -6843, 4208, 7199, -3599, -7504, 2964, 7753, -2312, -7949, 1643, 8086, -967, -8168, 283, 8190, 399, -8158, -1079, 8067, 1747, -7924, -2404, 7724, 3041, -7474, -3657, 7172, 4245, -6825, -4806, 6431, 5330, -5997, -5820, 5522, 6268, -5015, -6675, 4473, 7036, -3906, -7352, 3313, 7618, -2702, -7835, 2073, 8000, -1434, -8116, 787, 8177, -137, -8189, -513, 8148, 1156, -8057, -1793, 7915, 2414, -7727, -3021, 7489, 3606, -7208, -4169, 6883, 4704, -6518, -5211, 6113, 5683, -5675, -6122, 5202, 6521, -4702, -6883, 4173, 7202, -3624, -7479, 3053, 7711, -2468, -7899, 1868, 8040, -1261, -8136, 647, 8183, -33, -8187, -582, 8142, 1190, -8055, -1791, 7920, 2379, -7745, -2954, 7525, 3509, -7267, -4045, 6969, 4557, -6635, -5044, 6265, 5501, -5865, -5929, 5433, 6322, -4975, -6684, 4491, 7007, -3986, -7295, 3461, 7543, -2921, -7753, 2366, 7921, -1802, -8050, 1229, 8136, -654, -8183, 75, 8188, 501, -8153, -1074, 8077, 1639, -7964, -2196, 7810, 2738, -7620, -3268, 7393, 3778, -7133, -4271, 6838, 4740, -6514, -5187, 6158, 5607, -5776, -6001, 5367, 6365, -4937, -6700, 4483, 7002, -4012, -7272, 3523, 7508, -3021, -7711, 2506, 7877, -1983, -8009, 1451, 8104, -916, -8166, 377, 8190, 160, -8180, -696, 8134, 1226, -8055, -1751, 7940, 2265, -7795, -2770, 7615, 3259, -7406, -3736, 7166, 4193, -6899, -4634, 6603, 5053, -6283, -5452, 5937, 5826, -5571, -6178, 5182, 6502, -4776, -6802, 4350, 7072, -3911, -7315, 3457, 7528, -2993, -7714, 2517, 7868, -2035, -7993, 1545, 8087, -1054, -8152, 558, 8185, -63, -8189, -431, 8162, 921, -8108, -1408, 8023, 1885, -7912, -2357, 7771, 2816, -7605, -3266, 7412, 3701, -7196, -4124, 6953, 4529, -6690, -4919, 6404, 5290, -6099, -5643, 5772, 5974, -5430, -6287, 5069, 6575, -4695, -6843, 4305, 7087, -3905, -7308, 3492, 7504, -3071, -7677, 2641, 7824, -2205, -7947, 1763, 8044, -1319, -8118, 870, 8165, -423, -8189, -26, 8187, 472, -8162, -916, 8111, 1353, -8039, -1787, 7942, 2213, -7825, -2632, 7683, 3040, -7523, -3440, 7340, 3826, -7139, -4203, 6918, 4564, -6680, -4914, 6423, 5247, -6152, -5566, 5864, 5867, -5563, -6154, 5247, 6421, -4920, -6673, 4580, 6904, -4232, -7119, 3872, 7312, -3506, -7489, 3131, 7644, -2752, -7782, 2365, 7897, -1977, -7996, 1583, 8072, -1189, -8131, 792, 8169, -397, -8189, 1, 8188, 392, -8170, -784, 8132, 1170, -8077, -1554, 8003, 1931, -7913, -2304, 7804, 2669, -7680, -3027, 7538, 3376, -7383, -3718, 7211, 4048, -7026, -4371, 6826, 4680, -6614, -4981, 6388, 5268, -6152, -5546, 5903, 5808, -5645, -6060, 5375, 6297, -5098, -6523, 4810, 6733, -4516, -6931, 4214, 7113, -3907, -7283, 3592, 7436, -3274, -7577, 2949, 7702, -2623, -7814, 2292, 7910, -1960, -7993, 1625, 8060, -1290, -8114, 953, 8153, -618, -8179, 282, 8190, 51, -8189, -384, 8172, 713, -8144, -1041, 8102, 1364, -8048, -1684, 7981, 1999, -7903, -2310, 7811, 2615, -7710, -2916, 7596, 3208, -7474, -3497, 7338, 3777, -7195, -4051, 7041, 4317, -6879, -4576, 6706, 4826, -6527, -5070, 6338, 5304, -6144, -5530, 5940, 5747, -5731, -5956, 5514, 6154, -5294, -6345, 5065, 6525, -4834, -6698, 4596, 6859, -4355, -7013, 4109, 7155, -3861, -7290, 3608, 7414, -3355, -7530, 3097, 7634, -2839, -7731, 2577, 7817, -2316, -7895, 2052, 7962, -1790, -8022, 1525, 8071, -1263, -8113, 998, 8144, -737, -8169, 474, 8183, -215, -8191, -45, 8189, 301, -8180, -557, 8162, 809, -8138, -1060, 8104, 1307, -8066, -1553, 8018, 1793, -7965, -2033, 7903, 2266, -7837, -2498, 7763, 2725, -7684, -2949, 7598, 3168, -7508, -3384, 7410, 3593, -7309, -3801, 7202, 4001, -7091, -4200, 6974, 4391, -6854, -4580, 6728, 4762, -6600, -4941, 6466, 5113, -6331, -5282, 6191, 5444, -6049, -5603, 5902, 5754, -5755, -5903, 5603, 6045, -5450, -6184, 5293, 6316, -5137, -6444, 4976, 6566, -4816, -6684, 4653, 6796, -4490, -6905, 4324, 7007, -4159, -7106, 3991, 7198, -3824, -7288, 3655, 7371, -3488, -7451, 3318, 7525, -3151, -7596, 2981, 7661, -2813, -7724, 2644, 7780, -2477, -7834, 2309, 7882, -2143, -7928, 1976, 7969, -1812, -8007, 1646, 8040, -1484, -8071, 1321, 8096, -1161, -8120, 1000, 8139, -842, -8156, 684, 8168, -530, -8179, 375, 8185, -223, -8190, 71, 8190, 77, -8190, -225, 8185, 370, -8180, -514, 8170, 655, -8159, -796, 8145, 933, -8130, -1070, 8111, 1203, -8092, -1336, 8070, 1465, -8047, -1594, 8021, 1718, -7996, -1843, 7966, 1963, -7938, -2084, 7905, 2200, -7874, -2316, 7839, 2428, -7806, -2540, 7769, 2647, -7733, -2755, 7695, 2858, -7657, -2961, 7617, 3061, -7578, -3160, 7537, 3254, -7496, -3349, 7454, 3440, -7413, -3530, 7370, 3617, -7328, -3703, 7284, 3786, -7242, -3868, 7198, 3946, -7156, -4025, 7112, 4099, -7070, -4174, 7026, 4244, -6984, -4315, 6941, 4382, -6900, -4449, 6857, 4512, -6816, -4575, 6774, 4634, -6734, -4694, 6692, 4750, -6654, -4806, 6613, 4858, -6576, -4911, 6536, 4960, -6500, -5009, 6462, 5055, -6427, -5101, 6391, 5144, -6358, -5187, 6323, 5226, -6291, -5266, 6258, 5302, -6228, -5339, 6197, 5372, -6169, -5406, 6139, 5437, -6113, -5468, 6086, 5495, -6062, -5523, 6037, 5548, -6014, -5574, 5991, 5596, -5971, -5618, 5951, 5638, -5933, -5658, 5914, 5675, -5899, -5692, 5882, 5706, -5869, -5721, 5855, 5733, -5844, -5745, 5833, 5755, -5824, -5764, 5815, 5771, -5809, -5779, 5802, 5783, -5799, -5788, 5795, 5790, -5793, -5792, 5791, 5791, -5793, -5791, 5793, 5788, -5797, -5786, 5800, 5780, -5806, -5776, 5812, 5767, -5820, -5760, 5828, 5750, -5839, -5740, 5849, 5727, -5863, -5715, 5875, 5699, -5891, -5684, 5906, 5666, -5924, -5649, 5941, 5628, -5961, -5608, 5981, 5584, -6003, -5562, 6025, 5535, -6050, -5510, 6073, 5481, -6100, -5453, 6126, 5421, -6154, -5390, 6182, 5355, -6213, -5321, 6242, 5284, -6275, -5247, 6306, 5206, -6341, -5166, 6374, 5122, -6410, -5079, 6444, 5032, -6482, -4985, 6518, 4935, -6556, -4885, 6594, 4832, -6634, -4779, 6672, 4722, -6713, -4665, 6753, 4604, -6795, -4544, 6836, 4480, -6878, -4416, 6920, 4348, -6963, -4280, 7005, 4209, -7049, -4137, 7091, 4062, -7135, -3986, 7177, 3907, -7221, -3828, 7263, 3744, -7307, -3661, 7348, 3573, -7392, -3486, 7433, 3394, -7476, -3302, 7516, 3207, -7558, -3111, 7597, 3011, -7638, -2911, 7675, 2806, -7714, -2702, 7751, 2593, -7788, -2485, 7822, 2372, -7857, -2259, 7889, 2142, -7922, -2024, 7952, 1903, -7982, -1781, 8008, 1656, -8035, -1530, 8058, 1400, -8082, -1270, 8102, 1136, -8121, -1002, 8137, 864, -8153, -726, 8164, 584, -8175, -443, 8182, 297, -8188, -152, 8190, 2, -8191, 147, 8187, -299, -8183, 451, 8173, -607, -8163, 763, 8147, -921, -8130, 1080, 8108, -1241, -8084, 1402, 8055, -1565, -8024, 1728, 7988, -1894, -7949, 2059, 7905, -2226, -7859, 2392, 7807, -2561, -7753, 2728, 7692, -2898, -7630, 3065, 7561, -3235, -7489, 3403, 7411, -3572, -7330, 3739, 7243, -3908, -7153, 4074, 7057, -4242, -6957, 4406, 6851, -4572, -6741, 4734, 6625, -4897, -6506, 5056, 6380, -5216, -6251, 5372, 6115, -5527, -5975, 5678, 5829, -5829, -5680, 5975, 5523, -6121, -5364, 6261, 5197, -6400, -5028, 6533, 4851, -6665, -4672, 6791, 4486, -6915, -4296, 7032, 4101, -7147, -3902, 7256, 3697, -7361, -3490, 7459, 3276, -7554, -3059, 7641, 2837, -7725, -2613, 7800, 2382, -7872, -2150, 7934, 1913, -7993, -1674, 8042, 1430, -8086, -1185, 8122, 935, -8151, -684, 8172, 429, -8186, -174, 8190, -85, -8189, 344, 8177, -606, -8158, 867, 8129, -1131, -8094, 1393, 8047, -1658, -7994, 1921, 7929, -2185, -7857, 2446, 7774, -2708, -7684, 2967, 7582, -3226, -7473, 3481, 7353, -3736, -7225, 3985, 7085, -4233, -6938, 4476, 6779, -4716, -6613, 4950, 6436, -5181, -6252, 5404, 6056, -5624, -5853, 5836, 5639, -6043, -5419, 6241, 5187, -6434, -4950, 6617, 4702, -6794, -4448, 6960, 4184, -7120, -3915, 7268, 3637, -7408, -3354, 7536, 3062, -7655, -2766, 7762, 2463, -7859, -2156, 7943, 1842, -8017, -1525, 8076, 1202, -8125, -878, 8159, 548, -8183, -218, 8190, -116, -8187, 450, 8167, -786, -8136, 1121, 8088, -1458, -8029, 1792, 7953, -2127, -7864, 2457, 7759, -2787, -7642, 3112, 7508, -3434, -7362, 3749, 7199, -4061, -7024, 4365, 6833, -4665, -6630, 4954, 6411, -5238, -6181, 5510, 5936, -5775, -5679, 6028, 5408, -6272, -5127, 6502, 4832, -6722, -4527, 6927, 4210, -7121, -3885, 7298, 3548, -7463, -3203, 7611, 2848, -7744, -2488, 7860, 2118, -7960, -1744, 8042, 1363, -8107, -978, 8153, 588, -8182, -196, 8190, -199, -8182, 594, 8152, -991, -8105, 1386, 8036, -1780, -7950, 2171, 7841, -2559, -7716, 2941, 7568, -3320, -7403, 3689, 7217, -4053, -7014, 4406, 6790, -4752, -6550, 5084, 6289, -5407, -6013, 5714, 5718, -6010, -5409, 6289, 5082, -6554, -4741, 6801, 4385, -7031, -4017, 7242, 3634, -7434, -3242, 7605, 2837, -7757, -2424, 7886, 2000, -7994, -1572, 8078, 1135, -8140, -695, 8177, 249, -8191, 197, 8180, -647, -8145, 1094, 8084, -1542, -7999, 1984, 7888, -2424, -7754, 2856, 7593, -3283, -7410, 3699, 7200, -4107, -6968, 4501, 6712, -4884, -6434, 5251, 6133, -5604, -5812, 5937, 5468, -6254, -5107, 6549, 4726, -6825, -4329, 7077, 3914, -7307, -3486, 7511, 3042, -7692, -2588, 7844, 2122, -7971, -1648, 8069, 1164, -8139, -677, 8179, 184, -8191, 310, 8171, -806, -8124, 1299, 8043, -1791, -7935, 2276, 7794, -2756, -7625, 3226, 7425, -3686, -7198, 4132, 6940, -4565, -6656, 4980, 6343, -5379, -6006, 5756, 5642, -6114, -5256, 6446, 4846, -6755, -4417, 7035, 3966, -7290, -3500, 7514, 3016, -7709, -2519, 7871, 2009, -8002, -1490, 8098, 962, -8162, -429, 8189, -109, -8183, 646, 8139, -1184, -8062, 1717, 7947, -2246, -7799, 2765, 7613, -3274, -7395, 3769, 7141, -4251, -6855, 4712, 6536, -5155, -6187, 5575, 5807, -5971, -5401, 6339, 4966, -6680, -4509, 6989, 4027, -7268, -3526, 7511, 3004, -7720, -2469, 7891, 1918, -8026, -1358, 8120, 788, -8176, -214, 8190, -365, -8165, 941, 8098, -1517, -7991, 2085, 7841, -2645, -7653, 3192, 7423, -3726, -7156, 4240, 6850, -4736, -6508, 5206, 6129, -5653, -5719, 6068, 5275, -6455, -4804, 6806, 4304, -7123, -3780, 7401, 3233, -7641, -2669, 7837, 2086, -7993, -1492, 8104, 886, -8171, -276, 8190, -340, -8166, 954, 8093, -1566, -7976, 2169, 7810, -2763, -7601, 3340, 7345, -3902, -7048, 4440, 6707, -4956, -6327, 5442, 5906, -5899, -5452, 6320, 4961, -6706, -4441, 7050, 3890, -7355, -3317, 7613, 2719, -7828, -2106, 7992, 1475, -8109, -836, 8174, 188, -8190, 462, 8153, -1112, -8065, 1754, 7924, -2389, -7733, 3009, 7491, -3612, -7201, 4192, 6861, -4748, -6478, 5272, 6048, -5765, -5580, 6219, 5072, -6634, -4530, 7004, 3954, -7330, -3353, 7605, 2725, -7831, -2078, 8002, 1414, -8120, -741, 8181, 58, -8187, 624, 8133, -1306, -8025, 1979, 7858, -2641, -7636, 3284, 7358, -3907, -7028, 4502, 6645, -5068, -6215, 5596, 5736, -6087, -5217, 6532, 4656, -6933, -4061, 7281, 3433, -7578, -2780, 7818, 2102, -8001, -1409, 8122, 701, -8184, 11, 8182, -728, -8119, 1438, 7992, -2141, -7805, 2827, 7555, -3495, -7247, 4135, 6880, -4746, -6460, 5319, 5985, -5853, -5464, 6340, 4896, -6779, -4290, 7163, 3645, -7492, -2972, 7759, 2270, -7965, -1551, 8104, 815, -8179, -73, 8185, -674, -8125, 1415, 7994, -2147, -7798, 2862, 7535, -3555, -7208, 4219, 6818, -4849, -6371, 5438, 5866, -5983, -5311, 6476, 4707, -6916, -4063, 7294, 3380, -7612, -2667, 7861, 1928, -8043, -1171, 8153, 401, -8191, 373, 8155, -1147, -8047, 1910, 7865, -2660, -7612, 3385, 7288, -4083, -6898, 4743, 6442, -5363, -5927, 5932, 5354, -6450, -4733, 6906, 4063, -7301, -3356, 7626, 2614, -7881, -1847, 8060, 1059, -8165, -261, 8189, -543, -8137, 1341, 8004, -2131, -7795, 2899, 7508, -3642, -7148, 4350, 6715, -5018, -6218, 5635, 5655, -6200, -5037, 6703, 4365, -7141, -3650, 7506, 2895, -7799, -2111, 8010, 1302, -8143, -479, 8190, -351, -8156, 1178, 8035, -1997, -7832, 2794, 7546, -3566, -7182, 4301, 6741, -4993, -6229, 5632, 5648, -6215, -5009, 6731, 4312, -7178, -3570, 7547, 2786, -7837, -1972, 8042, 1134, -8161, -283, 8189, -575, -8130, 1426, 7979, -2265, -7742, 3078, 7417, -3861, -7011, 4601, 6523, -5292, -5963, 5924, 5333, -6492, -4644, 6985, 3898, -7402, -3109, 7733, 2280, -7978, -1426, 8130, 551, -8191, 329, 8154, -1210, -8025, 2076, 7799, -2921, -7483, 3732, 7077, -4502, -6588, 5219, 6018, -5877, -5377, 6463, 4669, -6976, -3905, 7403, 3091, -7744, -2240, 7990, 1357, -8141, -459, 8190, -449, -8142, 1351, 7991, -2240, -7743, 3101, 7396, -3927, -6959, 4703, 6432, -5424, -5825, 6077, 5141, -6655, -4394, 7149, 3587, -7555, -2735, 7863, 1845, -8073, -931, 8177, 1, -8178, 928, 8072, -1849, -7862, 2745, 7547, -3610, -7135, 4426, 6626, -5188, -6031, 5881, 5353, -6498, -4604, 7029, 3791, -7468, -2928, 7806, 2021, -8042, -1088, 8167, 136, -8184, 817, 8088, -1763, -7883, 2684, 7568, -3572, -7149, 4411, 6630, -5192, -6020, 5900, 5322, -6530, -4552, 7067, 3714, -7508, -2825, 7842, 1892, -8068, -933, 8178, -44, -8174, 1019, 8051, -1983, -7815, 2919, 7464, -3816, -7006, 4658, 6444, -5435, -5790, 6133, 5048, -6744, -4232, 7256, 3352, -7664, -2422, 7957, 1453, -8135, -463, 8190, -538, -8126, 1531, 7937, -2504, -7631, 3440, 7208, -4327, -6677, 5148, 6041, -5894, -5315, 6549, 4504, -7108, -3624, 7556, 2686, -7890, -1706, 8102, 696, -8189, 324, 8148, -1343, -7981, 2340, 7687, -3305, -7273, 4217, 6742, -5066, -6106, 5834, 5369, -6512, -4548, 7086, 3650, -7549, -2695, 7890, 1692, -8106, -663, 8189, -381, -8142, 1419, 7960, -2437, -7649, 3414, 7211, -4340, -6655, 5193, 5987, -5964, -5220, 6635, 4363, -7199, -3435, 7642, 2445, -7960, -1415, 8142, 358, -8190, 706, 8097, -1761, -7868, 2786, 7504, -3767, -7012, 4683, 6398, -5523, -5675, 6266, 4851, -6905, -3944, 7423, 2964, -7815, -1934, 8069, 866, -8185, 216, 8155, -1299, -7984, 2358, 7669, -3379, -7220, 4340, 6641, -5228, -5944, 6021, 5137, -6710, -4239, 7277, 3262, -7716, -2226, 8014, 1146, -8170, -45, 8175, -1059, -8033, 2145, 7741, -3194, -7309, 4185, 6740, -5102, -6047, 5924, 5240, -6639, -4335, 7229, 3346, -7688, -2296, 8001, 1198, -8166, -78, 8176, -1046, -8033, 2151, 7736, -3219, -7293, 4225, 6708, -5153, -5996, 5983, 5165, -6700, -4236, 7288, 3222, -7737, -2146, 8035, 1024, -8179, 117, 8161, -1260, -7986, 2377, 7652, -3452, -7168, 4458, 6540, -5379, -5784, 6193, 4909, -6887, -3938, 7443, 2884, -7852, -1773, 8102, 622, -8191, 541, 8113, -1696, -7873, 2817, 7470, -3884, -6916, 4872, 6218, -5763, -5394, 6535, 4455, -7176, -3426, 7667, 2322, -8002, -1170, 8170, -10, -8169, 1190, 7996, -2348, -7657, 3457, 7155, -4496, -6503, 5440, 5711, -6272, -4798, 6971, 3780, -7524, -2682, 7914, 1523, -8139, -332, 8186, -870, -8059, 2053, 7756, -3196, -7287, 4268, 6656, -5251, -5882, 6119, 4976, -6857, -3962, 7443, 2857, -7868, -1690, 8118, 481, -8190, 737, 8080, -1943, -7791, 3106, 7325, -4202, -6697, 5204, 5916, -6093, -5003, 6843, 3973, -7442, -2855, 7870, 1667, -8123, -442, 8189, -796, -8069, 2016, 7763, -3194, -7279, 4298, 6626, -5306, -5820, 6190, 4876, -6934, -3820, 7516, 2671, -7925, -1460, 8148, 211, -8181, 1042, 8020, -2275, -7671, 3453, 7139, -4554, -6438, 5545, 5582, -6408, -4593, 7117, 3490, -7658, -2305, 8015, 1061, -8180, 209, 8147, -1477, -7918, 2710, 7494, -3880, -6890, 4955, 6115, -5912, -5190, 6724, 4136, -7373, -2980, 7840, 1747, -8116, -471, 8189, -820, -8060, 2091, 7729, -3313, -7206, 4452, 6501, -5483, -5633, 6375, 4620, -7110, -3491, 7664, 2271, -8026, -993, 8183, -314, -8134, 1612, 7875, -2873, -7417, 4060, 6765, -5146, -5940, 6099, 4958, -6898, -3850, 7516, 2637, -7943, -1357, 8161, 38, -8168, 1283, 7959, -2573, -7543, 3795, 6926, -4921, -6128, 5916, 5164, -6758, -4064, 7419, 2853, -7886) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L32_i
    );

    L40_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (8040, 2216, -7678, -3471, 7111, 4630, -6357, -5667, 5434, 6550, -4369, -7261, 3188, 7778, -1926, -8092, 613, 8190, 713, -8076, -2021, 7748, 3273, -7220, -4440, 6503, 5488, -5619, -6394, 4588, 7132, -3441, -7686, 2204, 8040, -914, -8187, -400, 8122, 1700, -7851, -2958, 7377, 4137, -6717, -5211, 5884, 6149, -4904, -6931, 3799, 7535, -2601, -7950, 1336, 8161, -41, -8169, -1256, 7969, 2518, -7571, -3717, 6982, 4820, -6221, -5804, 5304, 6640, -4258, -7312, 3105, 7800, -1878, -8096, 605, 8190, 681, -8085, -1950, 7778, 3168, -7283, -4308, 6608, 5341, -5774, -6244, 4799, 6991, -3709, -7570, 2529, 7963, -1291, -8165, 21, 8167, 1246, -7975, -2484, 7589, 3659, -7023, -4747, 6288, 5718, -5406, -6554, 4393, 7230, -3280, -7737, 2087, 8057, -849, -8189, -410, 8125, 1657, -7871, -2864, 7432, 4002, -6820, -5046, 6048, 5969, -5137, -6754, 4105, 7379, -2982, -7835, 1788, 8106, -557, -8191, -688, 8086, 1914, -7796, -3097, 7327, 4205, -6691, -5218, 5902, 6108, -4981, -6861, 3945, 7454, -2823, -7880, 1637, 8126, -416, -8189, -814, 8066, 2022, -7764, -3186, 7286, 4275, -6648, -5270, 5860, 6144, -4944, -6882, 3918, 7464, -2807, -7883, 1634, 8125, -429, -8190, -787, 8072, 1982, -7779, -3135, 7315, 4215, -6693, -5204, 5924, 6077, -5029, -6819, 4024, 7410, -2935, -7843, 1782, 8104, -593, -8191, -608, 8101, 1793, -7840, -2941, 7409, 4022, -6823, -5019, 6090, 5905, -5231, -6668, 4260, 7286, -3202, -7752, 2076, 8053, -910, -8185, -276, 8144, 1453, -7935, -2601, 7559, 3691, -7028, -4704, 6349, 5618, -5542, -6415, 4619, 7078, -3604, -7596, 2514, 7955, -1376, -8153, 209, 8182, 959, -8046, -2108, 7744, 3211, -7288, -4250, 6682, 5199, -5944, -6044, 5086, 6765, -4128, -7350, 3086, 7786, -1986, -8068, 845, 8186, 309, -8143, -1458, 7937, 2574, -7576, -3640, 7064, 4631, -6415, -5532, 5639, 6321, -4755, -6987, 3777, 7514, -2729, -7895, 1626, 8121, -496, -8191, -645, 8101, 1770, -7856, -2861, 7458, 3894, -6919, -4854, 6247, 5717, -5457, -6471, 4563, 7100, -3585, -7595, 2538, 7943, -1446, -8143, 327, 8187, 796, -8079, -1904, 7817, 2973, -7412, -3987, 6866, 4924, -6195, -5769, 5408, 6505, -4523, -7121, 3554, 7603, -2523, -7947, 1444, 8141, -343, -8189, -766, 8084, 1857, -7835, -2915, 7440, 3917, -6914, -4849, 6261, 5689, -5497, -6428, 4634, 7049, -3690, -7544, 2680, 7901, -1625, -8119, 540, 8190, 551, -8118, -1633, 7900, 2683, -7544, -3686, 7054, 4621, -6442, -5475, 5716, 6231, -4894, -6878, 3984, 7403, -3009, -7801, 1980, 8061, -921, -8183, -155, 8161, 1225, -8002, -2275, 7703, 3282, -7274, -4234, 6720, 5110, -6055, -5901, 5285, 6588, -4429, -7165, 3497, 7618, -2509, -7944, 1478, 8135, -426, -8191, -634, 8108, 1680, -7892, -2698, 7544, 3669, -7073, -4579, 6483, 5411, -5790, -6154, 5000, 6794, -4131, -7323, 3194, 7731, -2208, -8013, 1185, 8163, -147, -8183, -895, 8068, 1919, -7826, -2912, 7456, 3856, -6969, -4738, 6369, 5542, -5670, -6258, 4880, 6872, -4016, -7378, 3088, 7765, -2113, -8031, 1105, 8169, -83, -8180, -941, 8062, 1946, -7820, -2923, 7455, 3850, -6976, -4719, 6389, 5512, -5706, -6220, 4934, 6831, -4089, -7337, 3181, 7729, -2228, -8005, 1240, 8157, -237, -8187, -771, 8091, 1763, -7876, -2730, 7541, 3652, -7095, -4521, 6541, 5319, -5893, -6038, 5157, 6665, -4347, -7195, 3471, 7615, -2548, -7925, 1587, 8117, -606, -8191, -385, 8143, 1367, -7980, -2329, 7698, 3254, -7308, -4133, 6811, 4950, -6218, -5696, 5535, 6357, -4776, -6929, 3948, 7399, -3066, -7765, 2141, 8019, -1188, -8161, 219, 8186, 751, -8098, -1711, 7895, 2643, -7584, -3539, 7165, 4383, -6650, -5167, 6041, 5876, -5352, -6505, 4588, 7042, -3764, -7483, 2888, 7820, -1976, -8051, 1036, 8171, -85, -8182, -867, 8080, 1804, -7872, -2718, 7556, 3592, -7142, -4418, 6630, 5183, -6034, -5879, 5355, 6495, -4609, -7025, 3802, 7461, -2947, -7799, 2053, 8033, -1136, -8164, 203, 8186, 730, -8104, -1653, 7915, 2552, -7626, -3418, 7238, 4238, -6759, -5003, 6192, 5702, -5549, -6329, 4835, 6873, -4062, -7331, 3237, 7693, -2375, -7961, 1482, 8126, -574, -8191, -342, 8152, 1250, -8013, -2144, 7774, 3007, -7440, -3835, 7014, 4611, -6504, -5332, 5913, 5985, -5253, -6566, 4528, 7064, -3751, -7477, 2928, 7798, -2073, -8027, 1192, 8156, -301, -8190, -595, 8124, 1480, -7964, -2349, 7707, 3186, -7362, -3987, 6928, 4737, -6416, -5432, 5828, 6061, -5174, -6621, 4459, 7100, -3696, -7499, 2889, 7808, -2052, -8029, 1190, 8156, -319, -8191, -557, 8130, 1423, -7979, -2274, 7737, 3096, -7409, -3883, 6996, 4623, -6507, -5313, 5945, 5940, -5319, -6502, 4633, 6989, -3898, -7399, 3120, 7726, -2311, -7969, 1475, 8123, -627, -8189, -228, 8164, 1078, -8053, -1917, 7853, 2732, -7570, -3518, 7205, 4263, -6765, -4963, 6252, 5607, -5674, -6192, 5036, 6709, -4348, -7157, 3612, 7526, -2842, -7818, 2042, 8026, -1224, -8151, 392, 8190, 440, -8147, -1269, 8017, 2081, -7807, -2872, 7515, 3631, -7150, -4354, 6710, 5029, -6205, -5653, 5636, 6218, -5013, -6722, 4339, 7155, -3624, -7518, 2873, 7804, -2096, -8013, 1298, 8141, -491, -8191, -322, 8158, 1128, -8048, -1924, 7857, 2698, -7592, -3447, 7252, 4159, -6844, -4831, 6370, 5454, -5837, -6026, 5247, 6537, -4611, -6987, 3930, 7369, -3214, -7682, 2468, 7920, -1702, -8086, 919, 8174, -131, -8187, -658, 8123, 1439, -7986, -2206, 7773, 2950, -7492, -3668, 7140, 4349, -6726, -4991, 6250, 5585, -5720, -6129, 5137, 6615, -4511, -7043, 3844, 7406, -3146, -7703, 2419, 7930, -1674, -8088, 914, 8173, -149, -8188, -618, 8129, 1376, -8002, -2123, 7803, 2848, -7539, -3550, 7209, 4217, -6820, -4849, 6370, 5437, -5869, -5979, 5318, 6467, -4724, -6902, 4090, 7276, -3424, -7591, 2729, 7839, -2014, -8024, 1282, 8139, -543, -8190, -201, 8171, 940, -8086, -1673, 7934, 2388, -7720, -3084, 7441, 3752, -7105, -4391, 6711, 4991, -6265, -5553, 5768, 6066, -5228, -6533, 4646, 6945, -4030, -7304, 3381, 7602, -2709, -7843, 2016, 8020, -1310, -8136, 593, 8187, 125, -8177, -842, 8102, 1550, -7968, -2247, 7771, 2923, -7518, -3578, 7206, 4202, -6842, -4796, 6426, 5351, -5965, -5866, 5459, 6335, -4914, -6759, 4333, 7130, -3723, -7449, 3085, 7712, -2428, -7920, 1752, 8068, -1067, -8160, 374, 8190, 319, -8164, -1010, 8078, 1690, -7937, -2359, 7737, 3008, -7486, -3637, 7180, 4237, -6827, -4808, 6425, 5342, -5981, -5841, 5495, 6296, -4974, -6709, 4418, 7073, -3835, -7390, 3225, 7655, -2597, -7869, 1950, 8028, -1293, -8135, 628, 8185, 39, -8183, -706, 8125, 1365, -8015, -2015, 7851, 2649, -7638, -3267, 7373, 3860, -7064, -4428, 6707, 4965, -6310, -5471, 5872, 5940, -5399, -6371, 4891, 6759, -4355, -7105, 3791, 7405, -3206, -7659, 2600, 7863, -1982, -8020, 1351, 8125, -714, -8182, 73, 8187, 565, -8144, -1201, 8049, 1826, -7908, -2440, 7718, 3037, -7485, -3616, 7205, 4170, -6884, -4701, 6522, 5200, -6125, -5670, 5690, 6104, -5225, -6503, 4729, 6862, -4209, -7182, 3663, 7459, -3100, -7694, 2518, 7883, -1926, -8029, 1321, 8127, -713, -8181, 100, 8188, 510, -8151, -1118, 8067, 1716, -7940, -2305, 7769, 2879, -7557, -3438, 7303, 3974, -7012, -4490, 6681, 4979, -6318, -5442, 5920, 5872, -5493, -6273, 5036, 6638, -4555, -6969, 4050, 7260, -3527, -7516, 2985, 7729, -2431, -7905, 1863, 8037, -1290, -8130, 709, 8180, -128, -8190, -455, 8157, 1031, -8085, -1604, 7971, 2164, -7819, -2715, 7628, 3249, -7401, -3768, 7137, 4265, -6840, -4743, 6509, 5194, -6150, -5621, 5760, 6018, -5345, -6388, 4904, 6724, -4443, -7030, 3960, 7300, -3462, -7538, 2947, 7738, -2422, -7903, 1884, 8030, -1342, -8122, 792, 8174, -243, -8191, -308, 8170, 855, -8114, -1398, 8019, 1932, -7892, -2458, 7727, 2970, -7531, -3469, 7301, 3950, -7042, -4415, 6751, 4857, -6433, -5279, 6087, 5676, -5717, -6049, 5323, 6394, -4909, -6714, 4473, 7002, -4022, -7262, 3553, 7490, -3073, -7688, 2580, 7852, -2079, -7986, 1569, 8085, -1057, -8153, 539, 8186, -22, -8188, -495, 8156, 1007, -8094, -1515, 7998, 2014, -7873, -2506, 7716, 2985, -7532, -3454, 7317, 3905, -7076, -4343, 6808, 4761, -6516, -5161, 6199, 5540, -5862, -5898, 5501, 6232, -5124, -6544, 4726, 6829, -4314, -7090, 3886, 7323, -3447, -7531, 2995, 7709, -2535, -7862, 2066, 7983, -1593, -8079, 1113, 8144, -633, -8182, 150, 8190, 330, -8172, -810, 8123, 1283, -8049, -1753, 7947, 2213, -7819, -2667, 7664, 3108, -7486, -3540, 7282, 3957, -7056, -4361, 6806, 4749, -6536, -5121, 6245, 5475, -5936, -5811, 5607, 6126, -5263, -6423, 4901, 6697, -4528, -6950, 4139, 7180, -3741, -7389, 3330, 7572, -2913, -7734, 2486, 7869, -2054, -7983, 1616, 8071, -1177, -8136, 733, 8175, -290, -8191, -154, 8182, 594, -8151, -1033, 8095, 1466, -8017, -1895, 7915, 2315, -7793, -2730, 7648, 3133, -7483, -3529, 7296, 3911, -7092, -4284, 6867, 4642, -6626, -4987, 6366, 5317, -6091, -5633, 5800, 5931, -5495, -6214, 5176, 6478, -4845, -6726, 4502, 6954, -4149, -7166, 3786, 7356, -3416, -7529, 3036, 7681, -2652, -7814, 2261, 7926, -1867, -8020, 1469, 8092, -1070, -8145, 667, 8177, -267, -8191, -135, 8184, 533, -8159, -930, 8113, 1322, -8050, -1711, 7966, 2093, -7867, -2471, 7748, 2840, -7613, -3203, 7460, 3556, -7293, -3902, 7108, 4235, -6910, -4560, 6696, 4872, -6469, -5174, 6228, 5462, -5976, -5739, 5710, 6001, -5435, -6252, 5148, 6486, -4853, -6708, 4547, 6913, -4235, -7106, 3913, 7281, -3587, -7443, 3253, 7587, -2915, -7718, 2571, 7831, -2225, -7931, 1875, 8012, -1524, -8080, 1169, 8130, -816, -8167, 460, 8186, -107, -8191, -247, 8180, 597, -8155, -947, 8114, 1291, -8060, -1634, 7990, 1971, -7907, -2305, 7810, 2631, -7701, -2953, 7577, 3267, -7442, -3576, 7293, 3876, -7135, -4170, 6963, 4454, -6782, -4731, 6589, 4997, -6388, -5256, 6175, 5504, -5955, -5743, 5725, 5970, -5488, -6189, 5242, 6395, -4990, -6593, 4730, 6777, -4466, -6953, 4195, 7115, -3920, -7267, 3638, 7407, -3354, -7536, 3065, 7652, -2774, -7759, 2479, 7852, -2184, -7935, 1884, 8005, -1586, -8065, 1284, 8112, -984, -8149, 683, 8173, -383, -8188, 83, 8190, 215, -8183, -512, 8164, 806, -8136, -1099, 8096, 1387, -8047, -1674, 7987, 1956, -7919, -2236, 7839, 2510, -7752, -2781, 7655, 3046, -7550, -3308, 7435, 3562, -7314, -3814, 7183, 4057, -7046, -4297, 6900, 4528, -6749, -4756, 6589, 4975, -6424, -5189, 6251, 5394, -6074, -5595, 5890, 5786, -5702, -5973, 5508, 6150, -5310, -6322, 5106, 6484, -4900, -6641, 4688, 6789, -4475, -6931, 4256, 7063, -4036, -7190, 3812, 7307, -3587, -7419, 3358, 7521, -3129, -7617, 2896, 7704, -2664, -7785, 2429, 7857, -2195, -7924, 1959, 7981, -1724, -8033, 1487, 8075, -1252, -8113, 1015, 8141, -781, -8165, 546, 8179, -313, -8189, 80, 8190, 150, -8187, -381, 8176, 608, -8160, -835, 8136, 1058, -8108, -1281, 8072, 1499, -8032, -1717, 7985, 1931, -7934, -2143, 7876, 2351, -7815, -2558, 7747, 2760, -7676, -2960, 7598, 3156, -7518, -3350, 7431, 3538, -7342, -3725, 7247, 3907, -7150, -4086, 7047, 4260, -6943, -4432, 6833, 4599, -6722, -4763, 6605, 4922, -6488, -5078, 6366, 5229, -6243, -5377, 6115, 5520, -5987, -5660, 5854, 5795, -5722, -5927, 5585, 6054, -5449, -6178, 5309, 6296, -5169, -6412, 5025, 6522, -4883, -6631, 4737, 6733, -4592, -6833, 4443, 6927, -4297, -7020, 4147, 7106, -3998, -7191, 3848, 7270, -3698, -7347, 3547, 7418, -3397, -7488, 3245, 7552, -3094, -7615, 2942, 7672, -2793, -7728, 2641, 7778, -2492, -7827, 2341, 7871, -2192, -7913, 2042, 7950, -1895, -7987, 1746, 8018, -1601, -8048, 1454, 8073, -1309, -8098, 1164, 8117, -1022, -8136, 879, 8150, -739, -8164, 598, 8173, -461, -8182, 322, 8187, -187, -8191, 51, 8190, 81, -8190, -214, 8186, 343, -8181, -473, 8173, 600, -8165, -727, 8152, 850, -8140, -974, 8125, 1095, -8110, -1215, 8091, 1332, -8072, -1450, 8051, 1564, -8030, -1678, 8005, 1788, -7981, -1899, 7954, 2006, -7928, -2113, 7899, 2217, -7871, -2320, 7840, 2421, -7810, -2521, 7777, 2618, -7745, -2715, 7711, 2808, -7678, -2901, 7642, 2991, -7608, -3081, 7571, 3168, -7536, -3255, 7498, 3338, -7462, -3421, 7423, 3501, -7387, -3581, 7348, 3657, -7310, -3734, 7271, 3807, -7234, -3880, 7194, 3950, -7156, -4021, 7117, 4087, -7079, -4154, 7040, 4218, -7002, -4282, 6963, 4343, -6926, -4404, 6887, 4461, -6851, -4519, 6813, 4574, -6777, -4629, 6739, 4681, -6704, -4733, 6667, 4782, -6633, -4832, 6597, 4878, -6563, -4925, 6528, 4968, -6496, -5012, 6462, 5053, -6431, -5094, 6398, 5133, -6368, -5172, 6337, 5207, -6308, -5244, 6278, 5277, -6251, -5311, 6222, 5342, -6196, -5374, 6169, 5402, -6145, -5431, 6119, 5458, -6096, -5485, 6072, 5509, -6051, -5533, 6029, 5555, -6009, -5578, 5989, 5597, -5971, -5618, 5952, 5635, -5936, -5653, 5919, 5669, -5905, -5685, 5890, 5698, -5878, -5712, 5864, 5723, -5854, -5736, 5843, 5745, -5834, -5755, 5825, 5762, -5818, -5770, 5811, 5775, -5806, -5781, 5800, 5785, -5798, -5789, 5794, 5790, -5793, -5792, 5791, 5791, -5793, -5792, 5793, 5789, -5796, -5787, 5798, 5783, -5803, -5779, 5808, 5772, -5815, -5767, 5821, 5758, -5830, -5750, 5838, 5740, -5849, -5730, 5859, 5717, -5871, -5706, 5883, 5691, -5898, -5677, 5912, 5661, -5928, -5645, 5944, 5626, -5962, -5608, 5979, 5587, -5999, -5567, 6018, 5544, -6040, -5522, 6061, 5496, -6085, -5472, 6107, 5444, -6132, -5417, 6156, 5388, -6183, -5358, 6208, 5326, -6237, -5295, 6264, 5260, -6293, -5226, 6322, 5189, -6353, -5153, 6382, 5113, -6415, -5074, 6446, 5032, -6479, -4991, 6512, 4946, -6546, -4902, 6579, 4854, -6615, -4808, 6649, 4757, -6686, -4708, 6721, 4655, -6758, -4602, 6794, 4546, -6832, -4491, 6869, 4432, -6907, -4374, 6944, 4312, -6983, -4251, 7021, 4186, -7060, -4122, 7098, 4054, -7137, -3986, 7175, 3915, -7214, -3844, 7252, 3770, -7291, -3696, 7329, 3619, -7368, -3541, 7405, 3460, -7443, -3380, 7479, 3296, -7517, -3212, 7553, 3124, -7590, -3037, 7625, 2946, -7661, -2855, 7694, 2761, -7729, -2667, 7761, 2569, -7794, -2471, 7825, 2370, -7856, -2269, 7885, 2165, -7914, -2060, 7941, 1952, -7969, -1844, 7993, 1733, -8018, -1621, 8040, 1506, -8062, -1392, 8081, 1274, -8101, -1156, 8117, 1034, -8133, -913, 8146, 788, -8159, -664, 8168, 536, -8178, -409, 8183, 278, -8189, -148, 8190, 14, -8191, 119, 8188, -255, -8185, 391, 8178, -530, -8170, 668, 8157, -809, -8144, 950, 8127, -1094, -8108, 1236, 8085, -1382, -8061, 1526, 8033, -1674, -8003, 1820, 7968, -1969, -7933, 2117, 7892, -2267, -7850, 2416, 7803, -2567, -7754, 2716, 7700, -2868, -7645, 3018, 7584, -3170, -7521, 3320, 7453, -3472, -7384, 3622, 7308, -3773, -7231, 3923, 7149, -4073, -7064, 4221, 6973, -4371, -6881, 4517, 6783, -4665, -6683, 4809, 6577, -4955, -6468, 5097, 6354, -5239, -6238, 5378, 6116, -5518, -5991, 5653, 5861, -5789, -5729, 5920, 5590, -6052, -5450, 6179, 5303, -6305, -5155, 6427, 5000, -6548, -4843, 6664, 4681, -6778, -4517, 6888, 4346, -6996, -4174, 7099, 3996, -7200, -3817, 7295, 3632, -7388, -3445, 7474, 3253, -7559, -3059, 7637, 2860, -7712, -2660, 7781, 2454, -7847, -2248, 7905, 2037, -7961, -1825, 8009, 1608, -8053, -1391, 8090, 1169, -8123, -947, 8148, 721, -8169, -495, 8182, 265, -8190, -36, 8190, -197, -8186, 429, 8172, -664, -8154, 897, 8127, -1134, -8095, 1369, 8054, -1606, -8008, 1841, 7953, -2078, -7892, 2312, 7822, -2547, -7746, 2780, 7661, -3013, -7571, 3243, 7470, -3473, -7365, 3699, 7249, -3925, -7128, 4146, 6998, -4366, -6861, 4582, 6716, -4795, -6564, 5003, 6404, -5209, -6237, 5409, 6062, -5606, -5881, 5796, 5691, -5983, -5496, 6163, 5292, -6339, -5083, 6507, 4865, -6670, -4643, 6825, 4413, -6974, -4178, 7115, 3936, -7250, -3689, 7375, 3435, -7494, -3178, 7603, 2914, -7705, -2646, 7796, 2373, -7881, -2097, 7953, 1815, -8019, -1532, 8072, 1243, -8118, -953, 8151, 659, -8176, -364, 8188, 66, -8191, 232, 8182, -533, -8163, 833, 8131, -1135, -8090, 1435, 8036, -1736, -7972, 2034, 7894, -2332, -7807, 2627, 7707, -2921, -7596, 3210, 7472, -3497, -7339, 3779, 7192, -4058, -7036, 4331, 6866, -4600, -6687, 4861, 6495, -5118, -6294, 5365, 6081, -5608, -5858, 5840, 5624, -6067, -5382, 6282, 5127, -6490, -4866, 6686, 4593, -6875, -4313, 7050, 4024, -7216, -3728, 7369, 3422, -7511, -3112, 7640, 2792, -7757, -2469, 7860, 2138, -7951, -1804, 8026, 1463, -8089, -1120, 8136, 772, -8170, -423, 8187, 70, -8191, 283, 8178, -638, -8151, 992, 8107, -1347, -8049, 1699, 7973, -2051, -7884, 2398, 7776, -2744, -7655, 3084, 7517, -3421, -7365, 3751, 7195, -4076, -7012, 4392, 6812, -4702, -6599, 5001, 6370, -5293, -6129, 5574, 5872, -5845, -5603, 6103, 5319, -6351, -5025, 6584, 4717, -6805, -4400, 7010, 4069, -7203, -3731, 7378, 3380, -7539, -3023, 7682, 2656, -7810, -2284, 7918, 1903, -8011, -1518, 8083, 1126, -8139, -732, 8173, 334, -8190, 65, 8186, -468, -8164, 868, 8120, -1270, -8059, 1668, 7975, -2065, -7873, 2457, 7749, -2845, -7608, 3226, 7445, -3602, -7264, 3968, 7062, -4327, -6843, 4674, 6604, -5012, -6349, 5337, 6074, -5650, -5784, 5947, 5476, -6231, -5154, 6497, 4816, -6749, -4465, 6981, 4099, -7197, -3722, 7392, 3332, -7568, -2933, 7722, 2523, -7857, -2106, 7968, 1680, -8059, -1250, 8125, 813, -8170, -375, 8189, -69, -8186, 511, 8158, -955, -8107, 1396, 8029, -1836, -7930, 2270, 7804, -2701, -7656, 3122, 7483, -3537, -7288, 3941, 7067, -4335, -6827, 4716, 6562, -5084, -6278, 5436, 5971, -5774, -5646, 6092, 5300, -6393, -4938, 6673, 4557, -6934, -4161, 7171, 3750, -7387, -3326, 7578, 2888, -7745, -2442, 7886, 1983, -8002, -1519, 8089, 1046, -8151, -571, 8184, 90, -8190, 391, 8166, -874, -8115, 1353, 8034, -1830, -7927, 2301, 7788, -2767, -7624, 3222, 7430, -3669, -7211, 4102, 6962, -4523, -6690, 4926, 6391, -5315, -6069, 5683, 5721, -6034, -5354, 6360, 4963, -6666, -4554, 6945, 4126, -7200, -3682, 7427, 3221, -7628, -2748, 7798, 2261, -7940, -1766, 8049, 1261, -8129, -752, 8176, 236, -8191, 280, 8173, -798, -8123, 1313, 8039, -1826, -7923, 2330, 7773, -2828, -7593, 3314, 7379, -3790, -7136, 4249, 6861, -4694, -6558, 5118, 6225, -5523, -5866, 5905, 5480, -6264, -5071, 6595, 4638, -6900, -4185, 7175, 3711, -7421, -3222, 7633, 2715, -7814, -2197, 7959, 1666, -8071, -1128, 8146, 582, -8186, -34, 8187, -518, -8153, 1067, 8080, -1614, -7972, 2154, 7824, -2686, -7643, 3206, 7423, -3714, -7170, 4204, 6881, -4677, -6561, 5127, 6206, -5556, -5824, 5958, 5410, -6334, -4972, 6678, 4506, -6993, -4020, 7273, 3510, -7519, -2985, 7728, 2441, -7900, -1886, 8032, 1318, -8126, -744, 8178, 163, -8191, 418, 8160, -1000, -8089, 1577, 7976, -2149, -7823, 2709, 7627, -3259, -7393, 3791, 7119, -4306, -6808, 4798, 6459, -5268, -6077, 5709, 5660, -6123, -5214, 6503, 4737, -6851, -4236, 7161, 3708, -7435, -3161, 7668, 2594, -7860, -2013, 8009, 1417, -8115, -815, 8175, 205, -8191, 406, 8159, -1018, -8084, 1624, 7961, -2224, -7795, 2810, 7581, -3384, -7326, 3938, 7027, -4472, -6688, 4980, 6308, -5462, -5892, 5911, 5439, -6329, -4955, 6708, 4438, -7050, -3897, 7349, 3328, -7608, -2741, 7819, 2134, -7985, -1515, 8102, 883, -8172, -247, 8190, -394, -8160, 1033, 8078, -1668, -7948, 2292, 7767, -2906, -7538, 3500, 7260, -4076, -6938, 4626, 6570, -5149, -6161, 5639, 5710, -6096, -5223, 6513, 4700, -6891, -4148, 7224, 3566, -7512, -2961, 7750, 2334, -7940, -1692, 8076, 1036, -8161, -373, 8190, -295, -8167, 961, 8088, -1623, -7956, 2275, 7768, -2914, -7530, 3533, 7237, -4131, -6897, 4700, 6508, -5240, -6074, 5743, 5596, -6209, -5080, 6631, 4526, -7010, -3941, 7339, 3325, -7619, -2687, 7843, 2026, -8015, -1352, 8128, 665, -8185, 27, 8182, -721, -8122, 1410, 8001, -2092, -7824, 2758, 7587, -3408, -7297, 4031, 6950, -4628, -6554, 5191, 6106, -5718, -5614, 6201, 5078, -6641, -4504, 7030, 3893, -7369, -3254, 7651, 2587, -7877, -1901, 8042, 1197, -8148, -485, 8190, -235, -8170, 952, 8085, -1665, -7939, 2364, 7730, -3049, -7461, 3708, 7131, -4342, -6746, 4941, 6306, -5504, -5816, 6022, 5277, -6495, -4697, 6914, 4076, -7281, -3422, 7588, 2738, -7836, -2033, 8018, 1307, -8137, -572, 8188, -172, -8173, 913, 8089, -1650, -7940, 2373, 7722, -3080, -7442, 3760, 7096, -4412, -6692, 5026, 6229, -5600, -5714, 6126, 5148, -6602, -4539, 7021, 3887, -7383, -3203, 7679, 2488, -7912, -1752, 8074, 998, -8168, -235, 8189, -532, -8140, 1295, 8018, -2050, -7826, 2785, 7562, -3500, -7233, 4182, 6836, -4830, -6380, 5434, 5863, -5992, -5294, 6495, 4675, -6941, -4014, 7324, 3312, -7642, -2582, 7888, 1824, -8064, -1050, 8164, 263, -8190, 525, 8139, -1313, -8013, 2087, 7810, -2845, -7535, 3576, 7186, -4276, -6771, 4934, 6289, -5549, -5747, 6110, 5148, -6615, -4501, 7056, 3807, -7431, -3077, 7733, 2314, -7962, -1529, 8112, 726, -8185, 84, 8176, -896, -8088, 1699, 7918, -2488, -7671, 3252, 7345, -3987, -6948, 4681, 6478, -5331, -5944, 5927, 5347, -6466, -4698, 6938, 3997, -7342, -3257, 7671, 2480, -7923, -1678, 8092, 856, -8180, -25, 8181, -809, -8100, 1634, 7932, -2446, -7683, 3231, 7351, -3986, -6943, 4697, 6459, -5363, -5908, 5970, 5291, -6517, -4619, 6994, 3895, -7398, -3129, 7721, 2327, -7964, -1500, 8119, 654, -8188, 199, 8166, -1053, -8057, 1895, 7858, -2719, -7574, 3513, 7204, -4272, -6755, 4982, 6229, -5640, -5635, 6234, 4975, -6762, -4260, 7212, 3494, -7584, -2689, 7869, 1851, -8067, -992, 8172, 119, -8185, 755, 8103, -1624, -7931, 2473, 7664, -3297, -7311, 4083, 6870, -4824, -6351, 5508, 5755, -6131, -5093, 6682, 4368, -7156, -3592, 7545, 2771, -7848, -1918, 8056, 1039, -8170, -148, 8185, -748, -8104, 1635, 7924, -2505, -7650, 3344, 7281, -4146, -6826, 4898, 6285, -5592, -5668, 6218, 4979, -6770, -4230, 7238, 3426, -7619, -2580, 7905, 1699, -8095, -798, 8183, -116, -8171, 1029, 8055, -1932, -7840, 2810, 7523, -3656, -7113, 4455, 6611, -5201, -6026, 5880, 5361, -6486, -4628, 7009, 3834, -7444, -2991, 7783, 2106, -8023, -1194, 8158, 264, -8189, 670, 8111, -1597, -7930, 2504, 7642, -3380, -7256, 4212, 6771, -4991, -6198, 5703, 5540, -6343, -4809, 6897, 4011, -7362, -3161, 7727, 2265, -7990, -1339, 8145, 391, -8191, 561, 8125, -1509, -7950, 2435, 7664, -3332, -7276, 4183, 6785, -4979, -6202, 5706, 5530, -6357, -4784, 6919, 3968, -7388, -3097, 7752, 2180, -8011, -1234, 8156, 266, -8189, 704, 8104, -1668, -7907, 2608, 7595, -3514, -7177, 4369, 6654, -5165, -6038, 5886, 5332, -6526, -4550, 7071, 3700, -7517, -2797, 7853, 1851, -8077, -878, 8181, -111, -8169, 1098, 8035, -2072, -7785, 3015, 7418, -3917, -6943, 4760, 6363, -5536, -5690, 6228, 4929, -6831, -4095, 7331, 3197, -7723, -2252, 7998, 1269, -8155, -268, 8187, -740, -8097, 1737, 7882, -2710, -7548, 3641, 7097, -4520, -6539, 5329, 5877, -6059, -5126, 6695, 4293, -7230, -3394, 7652, 2439, -7957, -1447, 8136, 429, -8191, 595, 8115, -1613, -7914, 2605, 7586, -3559, -7140, 4456, 6577, -5286, -5912, 6031, 5150, -6682, -4306, 7226, 3390, -7657, -2421, 7963, 1409, -8143, -376, 8189, -668, -8105, 1699, 7887, -2707, -7543, 3669, 7073, -4575, -6488, 5405, 5794, -6149, -5006, 6791, 4132, -7324, -3191, 7734, 2193, -8017, -1160, 8166, 104, -8180, 954, 8056, -1998, -7798, 3008, 7406, -3971, -6891, 4866, 6257, -5682, -5518, 6401, 4682, -7013, -3767, 7504, 2784, -7869, -1754, 8098, 691, -8190, 383, 8139, -1454, -7948, 2499, 7618, -3504, -7157, 4448, 6568, -5317, -5866, 6092, 5059, -6763, -4163, 7315, 3191, -7739, -2164, 8026, 1094, -8173, -6, 8173, -1085, -8029, 2156, 7740, -3193, -7313, 4171, 6753, -5078, -6073, 5892, 5280, -6603, -4393, 7193, 3424, -7655, -2392, 7977, 1314, -8156, -213, 8183, -896, -8063, 1988, 7792, -3046, -7380, 4048, 6829, -4978, -6152, 5814, 5359, -6546, -4466, 7155, 3488, -7633, -2445, 7966, 1353, -8153, -236, 8184, -889, -8063, 1996, 7787, -3069, -7366, 4083, 6801, -5022, -6109, 5865, 5297, -6599, -4385, 7205, 3386, -7676, -2322, 7997, 1210, -8166, -75, 8176, -1064, -8028, 2182, 7723, -3261, -7268, 4276, 6670, -5210, -5941, 6041, 5093, -6756, -4146, 7338, 3114, -7776, -2021, 8060, 885, -8186, 268, 8147, -1419, -7947, 2541, 7587, -3616, -7076, 4618, 6420, -5529, -5636, 6329, 4736, -7003, -3741, 7535, 2666, -7916, -1538, 8134, 376, -8189, 794, 8074, -1950, -7796, 3066, 7355, -4122, -6765, 5093, 6032, -5961, -5175, 6705, 4208, -7313, -3155, 7767, 2032, -8061, -868, 8186, -318, -8141, 1496, 7923, -2647, -7540, 3741, 6995, -4759, -6304, 5675, 5476, -6474, -4533, 7135, 3491, -7646, -2374, 7992, 1204, -8169, -8, 8169, -1191, -7995, 2364, 7647, -3489, -7135, 4538, 6465, -5492, -5657, 6325, 4722, -7023, -3686, 7567, 2565, -7948, -1389, 8153, 179, -8180, 1034, 8026, -2227, -7696, 3371, 7193, -4444, -6532, 5416, 5722, -6272, -4787, 6986, 3741, -7547, -2612, 7937, 1422, -8151, -200, 8180, -1030, -8026, 2236, 7689, -3394, -7179, 4475, 6503, -5457, -5680, 6314, 4725, -7029, -3662, 7583, 2512, -7965, -1306, 8162, 66, -8173, 1175, 7993, -2392, -7630, 3553, 7087, -4635, -6381, 5608, 5523, -6453, -4538, 7146, 3443, -7675, -2268, 8021, 1036, -8181, 219, 8146, -1473, -7921, 2691, 7505, -3848, -6913, 4914, 6154, -5865, -5249, 6675, 4215, -7329, -3081, 7805, 1870, -8096, -615, 8190, -658, -8089, 1915, 7790, -3129, -7304, 4266, 6637, -5303, -5811, 6209, 4839, -6967, -3750, 7553, 2566, -7956, -1320, 8162, 38, -8169, 1245, 7972, -2500, -7580, 3692, 6997, -4796, -6242, 5780, 5328, -6623, -4283, 7299, 3127, -7795, -1893, 8094, 609, -8191, 690, 8081, -1975, -7768, 3210, 7256, -4366, -6561, 5411, 5697, -6321, -4689, 7069, 3558, -7639, -2337, 8012, 1053, -8182, 257, 8139, -1565, -7889, 2831, 7433, -4028, -6786, 5119, 5960, -6081, -4981, 6883, 3869, -7509, -2656, 7937, 1371, -8160, -51, 8168, -1274, -7962, 2565, 7544, -3791, -6929, 4917, 6128, -5916, -5166, 6756, 4064, -7420, -2854, 7885) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L40_i
    );

process(Clk_96, Ce_F6 , TI , LG  )
    variable count: integer := 0;
    variable guard: boolean := False;
begin
    if TI = '1' then 	
	adress <= "11";
    elsif rising_edge(clk_96) then         
	    if LG = '0' and guard = False  then				 
		 guard := True;
		 adress <= adress +1;					 
		if adress = "11" then
		   adress <= "00";
		end if;
	    elsif LG = '1' then 
	       guard := False;
	    end if;	
    end if;					 
end process;

    pft_adress <= PFT & adress ;
process(PFT_adress, Rom_cos_L15_i, Rom_cos_L21_i, Rom_cos_L32_i, Rom_cos_L40_i)
begin
  if  pft_adress = "0110000000" or pft_adress = "0110001100" then
        Rom_cos_i <= Rom_cos_L15_i;
    elsif pft_adress = "0100000000" or pft_adress = "0100001100" then
        Rom_cos_i <= Rom_cos_L21_i;
    elsif pft_adress = "0010000000" or pft_adress = "0010001100" then
        Rom_cos_i <= Rom_cos_L32_i;
    elsif pft_adress = "0000000000" or pft_adress = "0000001100" or pft_adress = "1100000000" then
        Rom_cos_i <= Rom_cos_L40_i;
    end if; 
 end process;

process (Clk_96, Ce_F6, EN, Rom_cos_i )
begin
	 
    if EN = '1' then
       Rom_cos <= conv_std_logic_vector(Rom_cos_i- magic, data_rom);
    else
       Rom_cos <=(others => '0');
    end if;	
end process;end Behavioral;