
library IEEE;
        use IEEE.STD_LOGIC_1164.ALL;
        Use ieee.std_logic_arith.all;
        Use ieee.std_logic_unsigned.all;
        USE ieee.math_real.all;
        USE std.textio.ALL;
        USE IEEE.std_logic_textio.ALL;

library elementary;
        use elementary.s274types_pkg.all;
        use elementary.utility.all;
        use elementary.all;
    
entity MUX_signal_type3 is
       generic (
        
           data_pft: integer := 6;
                data_ppz : integer := 5;
                pft_widht : integer:= 6;
                pft_code : int_array := (10,27);
                data_rom : integer := 12
                                );
        Port(
                Clk_96 : in std_logic;
                Ce_F6 : in std_logic;
                En : in std_logic;      
                OD : in std_logic;              
                LG : in std_logic;              
                TI : in std_logic;
                PFT : in std_logic_vector (7 downto 0);         
                Sign_LCHM : in std_logic;
                Rom_cos : out std_logic_vector (13 downto 0)            
        );

end MUX_signal_type3;

architecture Behavioral of MUX_signal_type3 is

        signal P2_PFT : std_logic_vector(7 downto 0) := (others => '0');
    signal PFT_adress : std_logic_vector(9 downto 0) := (others => '0');
        signal Rom_cos_i : integer;
        signal adress : std_logic_vector(1 downto 0);  
        signal Rom_cos_L15_i : integer;
        signal Rom_cos_L15�31_i : integer;
        signal Rom_cos_L15�32_i : integer;
        signal Rom_cos_L15�33_i : integer;
        signal Rom_cos_L21_i : integer;
        signal Rom_cos_L21C31_i : integer;
        signal Rom_cos_L21C32_i : integer;
        signal Rom_cos_L21C33_i : integer;
        signal Rom_cos_L32_i : integer;
        signal Rom_cos_L32C31_i : integer;
        signal Rom_cos_L32C32_i : integer;
        signal Rom_cos_L32C33_i : integer;
begin

    L15_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-8146, -1520, 7899, 2795, -7449, -3996, 6805, 5089, -5990, -6049, 5021, 6851, -3930, -7478, 2739, 7912, -1485, -8148, 196, 8178, 1093, -8007, -2353, 7637, 3550, -7082, -4658, 6354, 5647, -5476, -6500, 4466, 7191, -3354, -7710, 2163, 8043, -927, -8186, -330, 8135, 1573, -7895, -2778, 7471, 3913, -6878, -4957, 6127, 5882, -5240, -6673, 4236, 7308, -3140, -7780, 1976, 8074, -773, -8190, -445, 8123, 1648, -7880, -2813, 7464, 3912, -6890, -4924, 6167, 5826, -5316, -6603, 4353, 7236, -3303, -7716, 2185, 8031, -1027, -8180, -151, 8157, 1320, -7969, -2461, 7617, 3545, -7113, -4557, 6466, 5472, -5693, -6277, 4808, 6952, -3832, -7491, 2782, 7879, -1683, -8114, 553, 8190, 582, -8111, -1704, 7875, 2788, -7493, -3818, 6968, 4770, -6317, -5633, 5549, 6387, -4683, -7022, 3732, 7526, -2719, -7893, 1657, 8114, -571, -8191, -523, 8121, 1602, -7909, -2651, 7557, 3649, -7077, -4582, 6474, 5430, -5764, -6185, 4956, 6830, -4068, -7359, 3113, 7761, -2112, -8034, 1077, 8172, -30, -8177, -1016, 8046, 2040, -7788, -3029, 7403, 3964, -6904, -4835, 6295, 5624, -5591, -6325, 4800, 6922, -3940, -7412, 3020, 7785, -2060, -8040, 1070, 8171, -69, -8180, -931, 8066, 1912, -7835, -2862, 7487, 3766, -7034, -4613, 6479, 5389, -5836, -6087, 5109, 6694, -4315, -7206, 3462, 7614, -2566, -7917, 1636, 8107, -689, -8189, -266, 8157, 1211, -8018, -2139, 7770, 3032, -7423, -3885, 6977, 4680, -6445, -5415, 5829, 6074, -5143, -6655, 4393, 7148, -3592, -7551, 2748, 7857, -1874, -8066, 980, 8173, -79, -8183, -821, 8092, 1706, -7907, -2569, 7626, 3396, -7260, -4181, 6808, 4913, -6281, -5587, 5683, 6193, -5024, -6728, 4310, 7183, -3552, -7558, 2757, 7846, -1936, -8050, 1096, 8163, -250, -8190, -597, 8127, 1432, -7981, -2250, 7750, 3039, -7442, -3796, 7057, 4508, -6603, -5173, 6083, 5782, -5506, -6332, 4876, 6814, -4202, -7231, 3488, 7573, -2747, -7842, 1980, 8034, -1200, -8152, 410, 8190, 377, -8155, -1160, 8043, 1926, -7861, -2673, 7607, 3391, -7288, -4077, 6905, 4723, -6465, -5325, 5970, 5878, -5427, -6379, 4840, 6822, -4216, -7208, 3559, 7531, -2877, -7792, 2174, 7986, -1458, -8118, 733, 8182, -7, -8184, -717, 8120, 1429, -7995, -2129, 7809, 2808, -7566, -3463, 7266, 4088, -6916, -4681, 6516, 5235, -6072, -5751, 5585, 6220, -5063, -6646, 4507, 7020, -3924, -7347, 3316, 7619, -2690, -7841, 2048, 8007, -1398, -8121, 741, 8180, -84, -8188, -572, 8141, 1218, -8046, -1855, 7899, 2475, -7706, -3078, 7465, 3657, -7183, -4213, 6857, 4738, -6496, -5235, 6096, 5696, -5666, -6125, 5205, 6514, -4719, -6867, 4208, 7177, -3679, -7449, 3132, 7677, -2573, -7865, 2002, 8009, -1426, -8112, 845, 8172, -265, -8191, -315, 8168, 887, -8107, -1454, 8005, 2007, -7868, -2550, 7692, 3075, -7483, -3584, 7240, 4072, -6967, -4540, 6663, 4982, -6333, -5402, 5976, 5793, -5598, -6159, 5197, 6495, -4779, -6803, 4342, 7079, -3893, -7327, 3429, 7542, -2957, -7728, 2475, 7880, -1989, -8004, 1497, 8094, -1005, -8156, 511, 8186, -21, -8188, -467, 8160, 948, -8105, -1424, 8021, 1890, -7912, -2347, 7777, 2792, -7618, -3225, 7435, 3643, -7231, -4049, 7005, 4436, -6761, -4809, 6497, 5162, -6218, -5499, 5920, 5816, -5611, -6115, 5286, 6393, -4952, -6653, 4604, 6890, -4250, -7110, 3886, 7306, -3516, -7485, 3139, 7641, -2760, -7778, 2376, 7894, -1991, -7992, 1603, 8068, -1217, -8127, 830, 8166, -447, -8188, 65, 8190, 312, -8176, -687, 8144, 1054, -8098, -1417, 8034, 1773, -7956, -2123, 7863, 2463, -7757, -2797, 7637, 3121, -7506, -3437, 7361, 3742, -7208, -4040, 7041, 4325, -6867, -4603, 6682, 4868, -6491, -5124, 6289, 5367, -6083, -5602, 5868, 5824, -5649, -6037, 5423, 6237, -5195, -6428, 4960, 6606, -4724, -6776, 4482, 6932, -4241, -7081, 3995, 7217, -3750, -7345, 3502, 7461, -3255, -7570, 3006, 7666, -2760, -7756, 2512, 7834, -2267, -7906, 2022, 7967, -1780, -8022, 1538, 8067, -1301, -8106, 1064, 8135, -832, -8160, 601, 8176, -375, -8187, 151, 8190, 68, -8190, -285, 8181, 496, -8169, -705, 8151, 908, -8129, -1109, 8101, 1303, -8071, -1495, 8035, 1680, -7997, -1863, 7954, 2040, -7910, -2213, 7862, 2381, -7812, -2545, 7759, 2703, -7705, -2858, 7647, 3007, -7590, -3153, 7530, 3292, -7470, -3429, 7407, 3560, -7346, -3688, 7282, 3810, -7220, -3929, 7155, 4042, -7093, -4153, 7028, 4257, -6966, -4360, 6903, 4456, -6842, -4551, 6780, 4639, -6721, -4726, 6661, 4807, -6603, -4886, 6546, 4960, -6491, -5032, 6436, 5098, -6385, -5163, 6334, 5223, -6286, -5281, 6238, 5334, -6194, -5386, 6150, 5433, -6110, -5478, 6070, 5519, -6035, -5559, 5999, 5593, -5968, -5627, 5938, 5656, -5912, -5684, 5886, 5707, -5865, -5730, 5844, 5748, -5828, -5765, 5812, 5777, -5801, -5789, 5791, 5796, -5785, -5802, 5780, 5804, -5779, -5805, 5779, 5802, -5784, -5798, 5789, 5789, -5799, -5780, 5810, 5766, -5825, -5751, 5841, 5732, -5861, -5712, 5882, 5687, -5907, -5661, 5933, 5631, -5963, -5600, 5994, 5563, -6029, -5526, 6064, 5484, -6104, -5441, 6143, 5393, -6187, -5344, 6231, 5289, -6278, -5233, 6326, 5172, -6377, -5110, 6428, 5042, -6483, -4972, 6537, 4897, -6594, -4821, 6651, 4738, -6711, -4654, 6770, 4564, -6832, -4472, 6893, 4375, -6956, -4275, 7018, 4169, -7083, -4061, 7145, 3946, -7210, -3830, 7272, 3707, -7336, -3581, 7397, 3450, -7460, -3315, 7520, 3175, -7581, -3031, 7638, 2881, -7696, -2729, 7750, 2570, -7804, -2408, 7854, 2240, -7903, -2069, 7947, 1891, -7991, -1711, 8029, 1524, -8066, -1335, 8096, 1139, -8125, -941, 8147, 737, -8167, -531, 8179, 318, -8189, -104, 8190, -116, -8188, 338, 8178, -566, -8163, 794, 8140, -1028, -8111, 1262, 8073, -1501, -8030, 1741, 7976, -1984, -7916, 2227, 7846, -2474, -7769, 2720, 7681, -2968, -7586, 3215, 7479, -3463, -7365, 3710, 7238, -3957, -7104, 4201, 6957, -4445, -6801, 4685, 6634, -4923, -6457, 5157, 6268, -5388, -6069, 5613, 5858, -5834, -5638, 6048, 5405, -6258, -5163, 6458, 4909, -6653, -4646, 6838, 4370, -7015, -4086, 7181, 3790, -7338, -3487, 7483, 3172, -7618, -2849, 7738, 2517, -7848, -2178, 7942, 1829, -8023, -1475, 8088, 1112, -8139, -746, 8171, 372, -8189, 4, 8188, -386, -8171, 769, 8134, -1156, -8080, 1541, 8005, -1929, -7912, 2314, 7797, -2699, -7665, 3079, 7510, -3457, -7337, 3827, 7141, -4192, -6927, 4548, 6691, -4897, -6437, 5233, 6160, -5560, -5866, 5872, 5550, -6171, -5218, 6453, 4866, -6720, -4497, 6967, 4111, -7197, -3710, 7404, 3292, -7591, -2863, 7753, 2418, -7893, -1964, 8005, 1498, -8094, -1025, 8153, 543, -8186, -58, 8188, -434, -8163, 926, 8106, -1420, -8020, 1910, 7902, -2399, -7754, 2880, 7574, -3355, -7364, 3819, 7121, -4272, -6849, 4709, 6546, -5132, -6215, 5535, 5853, -5918, -5466, 6277, 5051, -6613, -4612, 6919, 4148, -7199, -3664, 7446, 3157, -7662, -2635, 7841, 2095, -7987, -1543, 8093, 978, -8162, -407, 8190, -172, -8178, 752, 8124, -1334, -8029, 1910, 7890, -2483, -7711, 3043, 7488, -3593, -7224, 4125, 6918, -4639, -6574, 5129, 6189, -5595, -5768, 6030, 5310, -6434, -4820, 6802, 4298, -7134, -3748, 7423, 3171, -7670, -2573, 7871, 1954, -8026, -1321, 8129, 675, -8184, -22, 8185, -637, -8134, 1293, 8029, -1946, -7871, 2588, 7658, -3218, -7394, 3828, 7076, -4417, -6709, 4976, 6291, -5505, -5829, 5996, 5320, -6449, -4772, 6855, 4185, -7215, -3565, 7521, 2914, -7775, -2239, 7969, 1542, -8105, -831, 8177, 108, -8188, 617, 8132, -1343, -8012, 2060, 7826, -2767, -7577, 3452, 7263, -4114, -6889, 4742, 6453, -5337, -5962, 5886, 5416, -6390, -4823, 6839, 4182, -7232, -3504, 7560, 2789, -7825, -2048, 8019, 1283, -8142, -504, 8190, -285, -8163, 1073, 8058, -1857, -7878, 2625, 7621, -3373, -7290, 4090, 6885, -4772, -6413, 5408, 5873, -5996, -5274, 6524, 4618, -6990, -3913, 7385, 3163, -7707, -2378, 7949, 1564, -8110, -731, 8185, -115, -8174, 962, 8073, -1803, -7885, 2627, 7609, -3428, -7249, 4192, 6805, -4914, -6284, 5581, 5688, -6190, -5026, 6729, 4301, -7193, -3525, 7574, 2702, -7868, -1846, 8069, 963, -8175, -66, 8181, -837, -8090, 1732, 7897, -2611, -7607, 3459, 7219, -4269, -6740, 5027, 6172, -5725, -5525, 6351, 4802, -6899, -4016, 7357, 3172, -7722, -2284, 7984, 1361, -8143, -418, 8190, -536, -8129, 1485, 7954, -2419, -7670, 3322, 7277, -4183, -6783, 4987, 6189, -5725, -5507, 6382, 4741, -6952, -3906, 7422, 3009, -7787, -2067, 8036, 1088, -8170, -92, 8180, -911, -8069, 1903, 7834, -2870, -7480, 3796, 7008, -4668, -6427, 5469, 5742, -6189, -4967, 6813, 4108, -7332, -3182, 7734, 2200, -8014, -1181, 8164, 138, -8182, 910, 8064, -1949, -7814, 2956, 7431, -3920, -6923, 4819, 6294, -5641, -5558, 6368, 4722, -6989, -3804, 7489, 2814, -7862, -1773, 8096, 696, -8190, 396, 8136, -1486, -7938, 2551, 7594, -3575, -7112, 4536, 6496, -5418, -5761, 6201, 4915, -6874, -3975, 7417, 2956, -7825, -1880, 8083, 762, -8189, 372, 8136, -1505, -7928, 2609, 7562, -3669, -7049, 4658, 6392, -5559, -5609, 6351, 4709, -7020, -3713, 7547, 2637, -7924, -1506, 8138, 338, -8188, 839, 8066, -2003, -7777, 3128, 7323, -4192, -6714, 5169, 5959, -6040, -5076, 6783, 4080, -7384, -2994, 7824, 1837, -8097, -639, 8190, -579, -8105, 1786, 7838, -2958, -7396, 4066, 6784, -5087, -6019, 5994, 5112, -6769, -4088, 7388, 2964, -7840, -1770, 8109, 529, -8191, 726, 8078, -1969, -7776, 3167, 7286, -4296, -6621, 5322, 5793, -6224, -4824, 6976, 3733, -7561, -2549, 7960, 1297, -8165, -11, 8166, -1281, -7964, 2543, 7559, -3745, -6964, 4855, 6187, -5845, -5253, 6686, 4178, -7359, -2994, 7841, 1727, -8121, -413, 8187, -918, -8038, 2226, 7674, -3480, -7106, 4642, 6344, -5685, -5410)     
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L15_i
    );

    L15�31_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (8145, 1519, -7900, -2796, 7448, 3995, -6806, -5090, 5989, 6048, -5022, -6852, 3929, 7477, -2740, -7913, 1484, 8147, -197, -8179, -1094, 8006, 2352, -7638, -3551, 7081, 4657, -6355, -5648, 5475, 6499, -4467, -7192, 3353, 7709, -2164, -8044, 926, 8185, 329, -8136, -1574, 7894, 2777, -7472, -3914, 6877, 4956, -6128, -5883, 5239, 6672, -4237, -7309, 3139, 7779, -1977, -8075, 772, 8189, 444, -8124, -1649, 7879, 2812, -7465, -3913, 6889, 4923, -6168, -5827, 5315, 6602, -4354, -7237, 3302, 7715, -2186, -8032, 1026, 8179, 150, -8158, -1321, 7968, 2460, -7618, -3546, 7112, 4556, -6467, -5473, 5692, 6276, -4809, -6953, 3831, 7490, -2783, -7880, 1682, 8113, -554, -8191, -583, 8110, 1703, -7876, -2789, 7492, 3817, -6969, -4771, 6316, 5632, -5550, -6388, 4682, 7021, -3733, -7527, 2718, 7892, -1658, -8115, 570, 8190, 522, -8122, -1603, 7908, 2650, -7558, -3650, 7076, 4581, -6475, -5431, 5763, 6184, -4957, -6831, 4067, 7358, -3114, -7762, 2111, 8033, -1078, -8173, 29, 8176, 1015, -8047, -2041, 7787, 3028, -7404, -3965, 6903, 4834, -6296, -5625, 5590, 6324, -4801, -6923, 3939, 7411, -3021, -7786, 2059, 8039, -1071, -8172, 68, 8179, 930, -8067, -1913, 7834, 2861, -7488, -3767, 7033, 4612, -6480, -5390, 5835, 6086, -5110, -6695, 4314, 7205, -3463, -7615, 2565, 7916, -1637, -8108, 688, 8188, 265, -8158, -1212, 8017, 2138, -7771, -3033, 7422, 3884, -6978, -4681, 6444, 5414, -5830, -6075, 5142, 6654, -4394, -7149, 3591, 7550, -2749, -7858, 1873, 8065, -981, -8174, 78, 8182, 820, -8093, -1707, 7906, 2568, -7627, -3397, 7259, 4180, -6809, -4914, 6280, 5586, -5684, -6194, 5023, 6727, -4311, -7184, 3551, 7557, -2758, -7847, 1935, 8049, -1097, -8164, 249, 8189, 596, -8128, -1433, 7980, 2249, -7751, -3040, 7441, 3795, -7058, -4509, 6602, 5172, -6084, -5783, 5505, 6331, -4877, -6815, 4201, 7230, -3489, -7574, 2746, 7841, -1981, -8035, 1199, 8151, -411, -8191, -378, 8154, 1159, -8044, -1927, 7860, 2672, -7608, -3392, 7287, 4076, -6906, -4724, 6464, 5324, -5971, -5879, 5426, 6378, -4841, -6823, 4215, 7207, -3560, -7532, 2876, 7791, -2175, -7987, 1457, 8117, -734, -8183, 6, 8183, 716, -8121, -1430, 7994, 2128, -7810, -2809, 7565, 3462, -7267, -4089, 6915, 4680, -6517, -5236, 6071, 5750, -5586, -6221, 5062, 6645, -4508, -7021, 3923, 7346, -3317, -7620, 2689, 7840, -2049, -8008, 1397, 8120, -742, -8181, 83, 8187, 571, -8142, -1219, 8045, 1854, -7900, -2476, 7705, 3077, -7466, -3658, 7182, 4212, -6858, -4739, 6495, 5234, -6097, -5697, 5665, 6124, -5206, -6515, 4718, 6866, -4209, -7178, 3678, 7448, -3133, -7678, 2572, 7864, -2003, -8010, 1425, 8111, -846, -8173, 264, 8190, 314, -8169, -888, 8106, 1453, -8006, -2008, 7867, 2549, -7693, -3076, 7482, 3583, -7241, -4073, 6966, 4539, -6664, -4983, 6332, 5401, -5977, -5794, 5597, 6158, -5198, -6496, 4778, 6802, -4343, -7080, 3892, 7326, -3430, -7543, 2956, 7727, -2476, -7881, 1988, 8003, -1498, -8095, 1004, 8155, -512, -8187, 20, 8187, 466, -8161, -949, 8104, 1423, -8022, -1891, 7911, 2346, -7778, -2793, 7617, 3224, -7436, -3644, 7230, 4048, -7006, -4437, 6760, 4808, -6498, -5163, 6217, 5498, -5921, -5817, 5610, 6114, -5287, -6394, 4951, 6652, -4605, -6891, 4249, 7109, -3887, -7307, 3515, 7484, -3140, -7642, 2759, 7777, -2377, -7895, 1990, 7991, -1604, -8069, 1216, 8126, -831, -8167, 446, 8187, -66, -8191, -313, 8175, 686, -8145, -1055, 8097, 1416, -8035, -1774, 7955, 2122, -7864, -2464, 7756, 2796, -7638, -3122, 7505, 3436, -7362, -3743, 7207, 4039, -7042, -4326, 6866, 4602, -6683, -4869, 6490, 5123, -6290, -5368, 6082, 5601, -5869, -5825, 5648, 6036, -5424, -6238, 5194, 6427, -4961, -6607, 4723, 6775, -4483, -6933, 4240, 7080, -3996, -7218, 3749, 7344, -3503, -7462, 3254, 7569, -3007, -7667, 2759, 7755, -2513, -7835, 2266, 7905, -2023, -7968, 1779, 8021, -1539, -8068, 1300, 8105, -1065, -8136, 831, 8159, -602, -8177, 374, 8186, -152, -8191, -69, 8189, 284, -8182, -497, 8168, 704, -8152, -909, 8128, 1108, -8102, -1304, 8070, 1494, -8036, -1681, 7996, 1862, -7955, -2041, 7909, 2212, -7863, -2382, 7811, 2544, -7760, -2704, 7704, 2857, -7648, -3008, 7589, 3152, -7531, -3293, 7469, 3428, -7408, -3561, 7345, 3687, -7283, -3811, 7219, 3928, -7156, -4043, 7092, 4152, -7029, -4258, 6965, 4359, -6904, -4457, 6841, 4550, -6781, -4640, 6720, 4725, -6662, -4808, 6602, 4885, -6547, -4961, 6490, 5031, -6437, -5099, 6384, 5162, -6335, -5224, 6285, 5280, -6239, -5335, 6193, 5385, -6151, -5434, 6109, 5477, -6071, -5520, 6034, 5558, -6000, -5594, 5967, 5626, -5939, -5657, 5911, 5683, -5887, -5708, 5864, 5729, -5845, -5749, 5827, 5764, -5813, -5778, 5800, 5788, -5792, -5797, 5784, 5801, -5781, -5805, 5778, 5804, -5780, -5803, 5783, 5797, -5790, -5790, 5798, 5779, -5811, -5767, 5824, 5750, -5842, -5733, 5860, 5711, -5883, -5688, 5906, 5660, -5934, -5632, 5962, 5599, -5995, -5564, 6028, 5525, -6065, -5485, 6103, 5440, -6144, -5394, 6186, 5343, -6232, -5290, 6277, 5232, -6327, -5173, 6376, 5109, -6429, -5043, 6482, 4971, -6538, -4898, 6593, 4820, -6652, -4739, 6710, 4653, -6771, -4565, 6831, 4471, -6894, -4376, 6955, 4274, -7019, -4170, 7082, 4060, -7146, -3947, 7209, 3829, -7273, -3708, 7335, 3580, -7398, -3451, 7459, 3314, -7521, -3176, 7580, 3030, -7639, -2882, 7695, 2728, -7751, -2571, 7803, 2407, -7855, -2241, 7902, 2068, -7948, -1892, 7990, 1710, -8030, -1525, 8065, 1334, -8097, -1140, 8124, 940, -8148, -738, 8166, 530, -8180, -319, 8188, 103, -8191, 115, 8187, -339, -8179, 565, 8162, -795, -8141, 1027, 8110, -1263, -8074, 1500, 8029, -1742, -7977, 1983, 7915, -2228, -7847, 2473, 7768, -2721, -7682, 2967, 7585, -3216, -7480, 3462, 7364, -3711, -7239, 3956, 7103, -4202, -6958, 4444, 6800, -4686, -6635, 4922, 6456, -5158, -6269, 5387, 6068, -5614, -5859, 5833, 5637, -6049, -5406, 6257, 5162, -6459, -4910, 6652, 4645, -6839, -4371, 7014, 4085, -7182, -3791, 7337, 3486, -7484, -3173, 7617, 2848, -7739, -2518, 7847, 2177, -7943, -1830, 8022, 1474, -8089, -1113, 8138, 745, -8172, -373, 8188, -5, -8189, 385, 8170, -770, -8135, 1155, 8079, -1542, -8006, 1928, 7911, -2315, -7798, 2698, 7664, -3080, -7511, 3456, 7336, -3828, -7142, 4191, 6926, -4549, -6692, 4896, 6436, -5234, -6161, 5559, 5865, -5873, -5551, 6170, 5217, -6454, -4867, 6719, 4496, -6968, -4112, 7196, 3709, -7405, -3293, 7590, 2862, -7754, -2419, 7892, 1963, -8006, -1499, 8093, 1024, -8154, -544, 8185, 57, -8189, 433, 8162, -927, -8107, 1419, 8019, -1911, -7903, 2398, 7753, -2881, -7575, 3354, 7363, -3820, -7122, 4271, 6848, -4710, -6547, 5131, 6214, -5536, -5854, 5917, 5465, -6278, -5052, 6612, 4611, -6920, -4149, 7198, 3663, -7447, -3158, 7661, 2634, -7842, -2096, 7986, 1542, -8094, -979, 8161, 406, -8191, 171, 8177, -753, -8125, 1333, 8028, -1911, -7891, 2482, 7710, -3044, -7489, 3592, 7223, -4126, -6919, 4638, 6573, -5130, -6190, 5594, 5767, -6031, -5311, 6433, 4819, -6803, -4299, 7133, 3747, -7424, -3172, 7669, 2572, -7872, -1955, 8025, 1320, -8130, -676, 8183, 21, -8186, 636, 8133, -1294, -8030, 1945, 7870, -2589, -7659, 3217, 7393, -3829, -7077, 4416, 6708, -4977, -6292, 5504, 5828, -5997, -5321, 6448, 4771, -6856, -4186, 7214, 3564, -7522, -2915, 7774, 2238, -7970, -1543, 8104, 830, -8178, -109, 8187, -618, -8133, 1342, 8011, -2061, -7827, 2766, 7576, -3453, -7264, 4113, 6888, -4743, -6454, 5336, 5961, -5887, -5417, 6389, 4822, -6840, -4183, 7231, 3503, -7561, -2790, 7824, 2047, -8020, -1284, 8141, 503, -8191, 284, 8162, -1074, -8059, 1856, 7877, -2626, -7622, 3372, 7289, -4091, -6886, 4771, 6412, -5409, -5874, 5995, 5273, -6525, -4619, 6989, 3912, -7386, -3164, 7706, 2377, -7950, -1565, 8109, 730, -8186, 114, 8173, -963, -8074, 1802, 7884, -2628, -7610, 3427, 7248, -4193, -6806, 4913, 6283, -5582, -5689, 6189, 5025, -6730, -4302, 7192, 3524, -7575, -2703, 7867, 1845, -8070, -964, 8174, 65, -8182, 836, 8089, -1733, -7898, 2610, 7606, -3460, -7220, 4268, 6739, -5028, -6173, 5724, 5524, -6352, -4803, 6898, 4015, -7358, -3173, 7721, 2283, -7985, -1362, 8142, 417, -8191, 535, 8128, -1486, -7955, 2418, 7669, -3323, -7278, 4182, 6782, -4988, -6190, 5724, 5506, -6383, -4742, 6951, 3905, -7423, -3010, 7786, 2066, -8037, -1089, 8169, 91, -8181, 910, 8068, -1904, -7835, 2869, 7479, -3797, -7009, 4667, 6426, -5470, -5743, 6188, 4966, -6814, -4109, 7331, 3181, -7735, -2201, 8013, 1180, -8165, -139, 8181, -911, -8065, 1948, 7813, -2957, -7432, 3919, 6922, -4820, -6295, 5640, 5557, -6369, -4723, 6988, 3803, -7490, -2815, 7861, 1772, -8097, -697, 8189, -397, -8137, 1485, 7937, -2552, -7595, 3574, 7111, -4537, -6497, 5417, 5760, -6202, -4916, 6873, 3974, -7418, -2957, 7824, 1879, -8084, -763, 8188, -373, -8137, 1504, 7927, -2610, -7563, 3668, 7048, -4659, -6393, 5558, 5608, -6352, -4710, 7019, 3712, -7548, -2638, 7923, 1505, -8139, -339, 8187, -840, -8067, 2002, 7776, -3129, -7324, 4191, 6713, -5170, -5960, 6039, 5075, -6784, -4081, 7383, 2993, -7825, -1838, 8096, 638, -8191, 578, 8104, -1787, -7839, 2957, 7395, -4067, -6785, 5086, 6018, -5995, -5113, 6768, 4087, -7389, -2965, 7839, 1769, -8110, -530, 8190, -727, -8079, 1968, 7775, -3168, -7287, 4295, 6620, -5323, -5794, 6223, 4823, -6977, -3734, 7560, 2548, -7961, -1298, 8164, 10, -8167, 1280, 7963, -2544, -7560, 3744, 6963, -4856, -6188, 5844, 5252, -6687, -4179, 7358, 2993, -7842, -1728, 8120, 412, -8188, 917, 8037, -2227, -7675, 3479, 7105, -4643, -6345, 5684, 5409)    
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L15�31_i
    );

    L15�32_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-8146, -1520, 7899, 2795, -7449, -3996, 6805, 5089, -5990, -6049, 5021, 6851, -3930, -7478, 2739, 7912, -1485, -8148, 196, 8178, 1093, -8007, -2353, 7637, 3550, -7082, -4658, 6354, 5647, -5476, -6500, 4466, 7191, -3354, -7710, 2163, 8043, -927, -8186, -330, 8135, 1573, -7895, -2778, 7471, 3913, -6878, -4957, 6127, 5882, -5240, -6673, 4236, 7308, -3140, -7780, 1976, 8074, -773, -8190, -445, 8123, 1648, -7880, -2813, 7464, 3912, -6890, -4924, 6167, 5826, -5316, -6603, 4353, 7236, -3303, -7716, 2185, 8031, -1027, -8180, -151, 8157, 1320, -7969, -2461, 7617, 3545, -7113, -4557, 6466, 5472, -5693, -6277, 4808, 6952, -3832, -7491, 2782, 7879, -1683, -8114, 553, 8190, 582, -8111, -1704, 7875, 2788, -7493, -3818, 6968, 4770, -6317, -5633, 5549, 6387, -4683, -7022, 3732, 7526, -2719, -7893, 1657, 8114, -571, -8191, -523, 8121, 1602, -7909, -2651, 7557, 3649, -7077, -4582, 6474, 5430, -5764, -6185, 4956, 6830, -4068, -7359, 3113, 7761, -2112, -8034, 1077, 8172, -30, -8177, -1016, 8046, 2040, -7788, -3029, 7403, 3964, -6904, -4835, 6295, 5624, -5591, -6325, 4800, 6922, -3940, -7412, 3020, 7785, -2060, -8040, 1070, 8171, -69, -8180, -931, 8066, 1912, -7835, -2862, 7487, 3766, -7034, -4613, 6479, 5389, -5836, -6087, 5109, 6694, -4315, -7206, 3462, 7614, -2566, -7917, 1636, 8107, -689, -8189, -266, 8157, 1211, -8018, -2139, 7770, 3032, -7423, -3885, 6977, 4680, -6445, -5415, 5829, 6074, -5143, -6655, 4393, 7148, -3592, -7551, 2748, 7857, -1874, -8066, 980, 8173, -79, -8183, -821, 8092, 1706, -7907, -2569, 7626, 3396, -7260, -4181, 6808, 4913, -6281, -5587, 5683, 6193, -5024, -6728, 4310, 7183, -3552, -7558, 2757, 7846, -1936, -8050, 1096, 8163, -250, -8190, -597, 8127, 1432, -7981, -2250, 7750, 3039, -7442, -3796, 7057, 4508, -6603, -5173, 6083, 5782, -5506, -6332, 4876, 6814, -4202, -7231, 3488, 7573, -2747, -7842, 1980, 8034, -1200, -8152, 410, 8190, 377, -8155, -1160, 8043, 1926, -7861, -2673, 7607, 3391, -7288, -4077, 6905, 4723, -6465, -5325, 5970, 5878, -5427, -6379, 4840, 6822, -4216, -7208, 3559, 7531, -2877, -7792, 2174, 7986, -1458, -8118, 733, 8182, -7, -8184, -717, 8120, 1429, -7995, -2129, 7809, 2808, -7566, -3463, 7266, 4088, -6916, -4681, 6516, 5235, -6072, -5751, 5585, 6220, -5063, -6646, 4507, 7020, -3924, -7347, 3316, 7619, -2690, -7841, 2048, 8007, -1398, -8121, 741, 8180, -84, -8188, -572, 8141, 1218, -8046, -1855, 7899, 2475, -7706, -3078, 7465, 3657, -7183, -4213, 6857, 4738, -6496, -5235, 6096, 5696, -5666, -6125, 5205, 6514, -4719, -6867, 4208, 7177, -3679, -7449, 3132, 7677, -2573, -7865, 2002, 8009, -1426, -8112, 845, 8172, -265, -8191, -315, 8168, 887, -8107, -1454, 8005, 2007, -7868, -2550, 7692, 3075, -7483, -3584, 7240, 4072, -6967, -4540, 6663, 4982, -6333, -5402, 5976, 5793, -5598, -6159, 5197, 6495, -4779, -6803, 4342, 7079, -3893, -7327, 3429, 7542, -2957, -7728, 2475, 7880, -1989, -8004, 1497, 8094, -1005, -8156, 511, 8186, -21, -8188, -467, 8160, 948, -8105, -1424, 8021, 1890, -7912, -2347, 7777, 2792, -7618, -3225, 7435, 3643, -7231, -4049, 7005, 4436, -6761, -4809, 6497, 5162, -6218, -5499, 5920, 5816, -5611, -6115, 5286, 6393, -4952, -6653, 4604, 6890, -4250, -7110, 3886, 7306, -3516, -7485, 3139, 7641, -2760, -7778, 2376, 7894, -1991, -7992, 1603, 8068, -1217, -8127, 830, 8166, -447, -8188, 65, 8190, 312, -8176, -687, 8144, 1054, -8098, -1417, 8034, 1773, -7956, -2123, 7863, 2463, -7757, -2797, 7637, 3121, -7506, -3437, 7361, 3742, -7208, -4040, 7041, 4325, -6867, -4603, 6682, 4868, -6491, -5124, 6289, 5367, -6083, -5602, 5868, 5824, -5649, -6037, 5423, 6237, -5195, -6428, 4960, 6606, -4724, -6776, 4482, 6932, -4241, -7081, 3995, 7217, -3750, -7345, 3502, 7461, -3255, -7570, 3006, 7666, -2760, -7756, 2512, 7834, -2267, -7906, 2022, 7967, -1780, -8022, 1538, 8067, -1301, -8106, 1064, 8135, -832, -8160, 601, 8176, -375, -8187, 151, 8190, 68, -8190, -285, 8181, 496, -8169, -705, 8151, 908, -8129, -1109, 8101, 1303, -8071, -1495, 8035, 1680, -7997, -1863, 7954, 2040, -7910, -2213, 7862, 2381, -7812, -2545, 7759, 2703, -7705, -2858, 7647, 3007, -7590, -3153, 7530, 3292, -7470, -3429, 7407, 3560, -7346, -3688, 7282, 3810, -7220, -3929, 7155, 4042, -7093, -4153, 7028, 4257, -6966, -4360, 6903, 4456, -6842, -4551, 6780, 4639, -6721, -4726, 6661, 4807, -6603, -4886, 6546, 4960, -6491, -5032, 6436, 5098, -6385, -5163, 6334, 5223, -6286, -5281, 6238, 5334, -6194, -5386, 6150, 5433, -6110, -5478, 6070, 5519, -6035, -5559, 5999, 5593, -5968, -5627, 5938, 5656, -5912, -5684, 5886, 5707, -5865, -5730, 5844, 5748, -5828, -5765, 5812, 5777, -5801, -5789, 5791, 5796, -5785, -5802, 5780, 5804, -5779, -5805, 5779, 5802, -5784, -5798, 5789, 5789, -5799, -5780, 5810, 5766, -5825, -5751, 5841, 5732, -5861, -5712, 5882, 5687, -5907, -5661, 5933, 5631, -5963, -5600, 5994, 5563, -6029, -5526, 6064, 5484, -6104, -5441, 6143, 5393, -6187, -5344, 6231, 5289, -6278, -5233, 6326, 5172, -6377, -5110, 6428, 5042, -6483, -4972, 6537, 4897, -6594, -4821, 6651, 4738, -6711, -4654, 6770, 4564, -6832, -4472, 6893, 4375, -6956, -4275, 7018, 4169, -7083, -4061, 7145, 3946, -7210, -3830, 7272, 3707, -7336, -3581, 7397, 3450, -7460, -3315, 7520, 3175, -7581, -3031, 7638, 2881, -7696, -2729, 7750, 2570, -7804, -2408, 7854, 2240, -7903, -2069, 7947, 1891, -7991, -1711, 8029, 1524, -8066, -1335, 8096, 1139, -8125, -941, 8147, 737, -8167, -531, 8179, 318, -8189, -104, 8190, -116, -8188, 338, 8178, -566, -8163, 794, 8140, -1028, -8111, 1262, 8073, -1501, -8030, 1741, 7976, -1984, -7916, 2227, 7846, -2474, -7769, 2720, 7681, -2968, -7586, 3215, 7479, -3463, -7365, 3710, 7238, -3957, -7104, 4201, 6957, -4445, -6801, 4685, 6634, -4923, -6457, 5157, 6268, -5388, -6069, 5613, 5858, -5834, -5638, 6048, 5405, -6258, -5163, 6458, 4909, -6653, -4646, 6838, 4370, -7015, -4086, 7181, 3790, -7338, -3487, 7483, 3172, -7618, -2849, 7738, 2517, -7848, -2178, 7942, 1829, -8023, -1475, 8088, 1112, -8139, -746, 8171, 372, -8189, 4, 8188, -386, -8171, 769, 8134, -1156, -8080, 1541, 8005, -1929, -7912, 2314, 7797, -2699, -7665, 3079, 7510, -3457, -7337, 3827, 7141, -4192, -6927, 4548, 6691, -4897, -6437, 5233, 6160, -5560, -5866, 5872, 5550, -6171, -5218, 6453, 4866, -6720, -4497, 6967, 4111, -7197, -3710, 7404, 3292, -7591, -2863, 7753, 2418, -7893, -1964, 8005, 1498, -8094, -1025, 8153, 543, -8186, -58, 8188, -434, -8163, 926, 8106, -1420, -8020, 1910, 7902, -2399, -7754, 2880, 7574, -3355, -7364, 3819, 7121, -4272, -6849, 4709, 6546, -5132, -6215, 5535, 5853, -5918, -5466, 6277, 5051, -6613, -4612, 6919, 4148, -7199, -3664, 7446, 3157, -7662, -2635, 7841, 2095, -7987, -1543, 8093, 978, -8162, -407, 8190, -172, -8178, 752, 8124, -1334, -8029, 1910, 7890, -2483, -7711, 3043, 7488, -3593, -7224, 4125, 6918, -4639, -6574, 5129, 6189, -5595, -5768, 6030, 5310, -6434, -4820, 6802, 4298, -7134, -3748, 7423, 3171, -7670, -2573, 7871, 1954, -8026, -1321, 8129, 675, -8184, -22, 8185, -637, -8134, 1293, 8029, -1946, -7871, 2588, 7658, -3218, -7394, 3828, 7076, -4417, -6709, 4976, 6291, -5505, -5829, 5996, 5320, -6449, -4772, 6855, 4185, -7215, -3565, 7521, 2914, -7775, -2239, 7969, 1542, -8105, -831, 8177, 108, -8188, 617, 8132, -1343, -8012, 2060, 7826, -2767, -7577, 3452, 7263, -4114, -6889, 4742, 6453, -5337, -5962, 5886, 5416, -6390, -4823, 6839, 4182, -7232, -3504, 7560, 2789, -7825, -2048, 8019, 1283, -8142, -504, 8190, -285, -8163, 1073, 8058, -1857, -7878, 2625, 7621, -3373, -7290, 4090, 6885, -4772, -6413, 5408, 5873, -5996, -5274, 6524, 4618, -6990, -3913, 7385, 3163, -7707, -2378, 7949, 1564, -8110, -731, 8185, -115, -8174, 962, 8073, -1803, -7885, 2627, 7609, -3428, -7249, 4192, 6805, -4914, -6284, 5581, 5688, -6190, -5026, 6729, 4301, -7193, -3525, 7574, 2702, -7868, -1846, 8069, 963, -8175, -66, 8181, -837, -8090, 1732, 7897, -2611, -7607, 3459, 7219, -4269, -6740, 5027, 6172, -5725, -5525, 6351, 4802, -6899, -4016, 7357, 3172, -7722, -2284, 7984, 1361, -8143, -418, 8190, -536, -8129, 1485, 7954, -2419, -7670, 3322, 7277, -4183, -6783, 4987, 6189, -5725, -5507, 6382, 4741, -6952, -3906, 7422, 3009, -7787, -2067, 8036, 1088, -8170, -92, 8180, -911, -8069, 1903, 7834, -2870, -7480, 3796, 7008, -4668, -6427, 5469, 5742, -6189, -4967, 6813, 4108, -7332, -3182, 7734, 2200, -8014, -1181, 8164, 138, -8182, 910, 8064, -1949, -7814, 2956, 7431, -3920, -6923, 4819, 6294, -5641, -5558, 6368, 4722, -6989, -3804, 7489, 2814, -7862, -1773, 8096, 696, -8190, 396, 8136, -1486, -7938, 2551, 7594, -3575, -7112, 4536, 6496, -5418, -5761, 6201, 4915, -6874, -3975, 7417, 2956, -7825, -1880, 8083, 762, -8189, 372, 8136, -1505, -7928, 2609, 7562, -3669, -7049, 4658, 6392, -5559, -5609, 6351, 4709, -7020, -3713, 7547, 2637, -7924, -1506, 8138, 338, -8188, 839, 8066, -2003, -7777, 3128, 7323, -4192, -6714, 5169, 5959, -6040, -5076, 6783, 4080, -7384, -2994, 7824, 1837, -8097, -639, 8190, -579, -8105, 1786, 7838, -2958, -7396, 4066, 6784, -5087, -6019, 5994, 5112, -6769, -4088, 7388, 2964, -7840, -1770, 8109, 529, -8191, 726, 8078, -1969, -7776, 3167, 7286, -4296, -6621, 5322, 5793, -6224, -4824, 6976, 3733, -7561, -2549, 7960, 1297, -8165, -11, 8166, -1281, -7964, 2543, 7559, -3745, -6964, 4855, 6187, -5845, -5253, 6686, 4178, -7359, -2994, 7841, 1727, -8121, -413, 8187, -918, -8038, 2226, 7674, -3480, -7106, 4642, 6344, -5685, -5410)     
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L15�32_i
    );

    L15�33_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (8145, 1519, -7900, -2796, 7448, 3995, -6806, -5090, 5989, 6048, -5022, -6852, 3929, 7477, -2740, -7913, 1484, 8147, -197, -8179, -1094, 8006, 2352, -7638, -3551, 7081, 4657, -6355, -5648, 5475, 6499, -4467, -7192, 3353, 7709, -2164, -8044, 926, 8185, 329, -8136, -1574, 7894, 2777, -7472, -3914, 6877, 4956, -6128, -5883, 5239, 6672, -4237, -7309, 3139, 7779, -1977, -8075, 772, 8189, 444, -8124, -1649, 7879, 2812, -7465, -3913, 6889, 4923, -6168, -5827, 5315, 6602, -4354, -7237, 3302, 7715, -2186, -8032, 1026, 8179, 150, -8158, -1321, 7968, 2460, -7618, -3546, 7112, 4556, -6467, -5473, 5692, 6276, -4809, -6953, 3831, 7490, -2783, -7880, 1682, 8113, -554, -8191, -583, 8110, 1703, -7876, -2789, 7492, 3817, -6969, -4771, 6316, 5632, -5550, -6388, 4682, 7021, -3733, -7527, 2718, 7892, -1658, -8115, 570, 8190, 522, -8122, -1603, 7908, 2650, -7558, -3650, 7076, 4581, -6475, -5431, 5763, 6184, -4957, -6831, 4067, 7358, -3114, -7762, 2111, 8033, -1078, -8173, 29, 8176, 1015, -8047, -2041, 7787, 3028, -7404, -3965, 6903, 4834, -6296, -5625, 5590, 6324, -4801, -6923, 3939, 7411, -3021, -7786, 2059, 8039, -1071, -8172, 68, 8179, 930, -8067, -1913, 7834, 2861, -7488, -3767, 7033, 4612, -6480, -5390, 5835, 6086, -5110, -6695, 4314, 7205, -3463, -7615, 2565, 7916, -1637, -8108, 688, 8188, 265, -8158, -1212, 8017, 2138, -7771, -3033, 7422, 3884, -6978, -4681, 6444, 5414, -5830, -6075, 5142, 6654, -4394, -7149, 3591, 7550, -2749, -7858, 1873, 8065, -981, -8174, 78, 8182, 820, -8093, -1707, 7906, 2568, -7627, -3397, 7259, 4180, -6809, -4914, 6280, 5586, -5684, -6194, 5023, 6727, -4311, -7184, 3551, 7557, -2758, -7847, 1935, 8049, -1097, -8164, 249, 8189, 596, -8128, -1433, 7980, 2249, -7751, -3040, 7441, 3795, -7058, -4509, 6602, 5172, -6084, -5783, 5505, 6331, -4877, -6815, 4201, 7230, -3489, -7574, 2746, 7841, -1981, -8035, 1199, 8151, -411, -8191, -378, 8154, 1159, -8044, -1927, 7860, 2672, -7608, -3392, 7287, 4076, -6906, -4724, 6464, 5324, -5971, -5879, 5426, 6378, -4841, -6823, 4215, 7207, -3560, -7532, 2876, 7791, -2175, -7987, 1457, 8117, -734, -8183, 6, 8183, 716, -8121, -1430, 7994, 2128, -7810, -2809, 7565, 3462, -7267, -4089, 6915, 4680, -6517, -5236, 6071, 5750, -5586, -6221, 5062, 6645, -4508, -7021, 3923, 7346, -3317, -7620, 2689, 7840, -2049, -8008, 1397, 8120, -742, -8181, 83, 8187, 571, -8142, -1219, 8045, 1854, -7900, -2476, 7705, 3077, -7466, -3658, 7182, 4212, -6858, -4739, 6495, 5234, -6097, -5697, 5665, 6124, -5206, -6515, 4718, 6866, -4209, -7178, 3678, 7448, -3133, -7678, 2572, 7864, -2003, -8010, 1425, 8111, -846, -8173, 264, 8190, 314, -8169, -888, 8106, 1453, -8006, -2008, 7867, 2549, -7693, -3076, 7482, 3583, -7241, -4073, 6966, 4539, -6664, -4983, 6332, 5401, -5977, -5794, 5597, 6158, -5198, -6496, 4778, 6802, -4343, -7080, 3892, 7326, -3430, -7543, 2956, 7727, -2476, -7881, 1988, 8003, -1498, -8095, 1004, 8155, -512, -8187, 20, 8187, 466, -8161, -949, 8104, 1423, -8022, -1891, 7911, 2346, -7778, -2793, 7617, 3224, -7436, -3644, 7230, 4048, -7006, -4437, 6760, 4808, -6498, -5163, 6217, 5498, -5921, -5817, 5610, 6114, -5287, -6394, 4951, 6652, -4605, -6891, 4249, 7109, -3887, -7307, 3515, 7484, -3140, -7642, 2759, 7777, -2377, -7895, 1990, 7991, -1604, -8069, 1216, 8126, -831, -8167, 446, 8187, -66, -8191, -313, 8175, 686, -8145, -1055, 8097, 1416, -8035, -1774, 7955, 2122, -7864, -2464, 7756, 2796, -7638, -3122, 7505, 3436, -7362, -3743, 7207, 4039, -7042, -4326, 6866, 4602, -6683, -4869, 6490, 5123, -6290, -5368, 6082, 5601, -5869, -5825, 5648, 6036, -5424, -6238, 5194, 6427, -4961, -6607, 4723, 6775, -4483, -6933, 4240, 7080, -3996, -7218, 3749, 7344, -3503, -7462, 3254, 7569, -3007, -7667, 2759, 7755, -2513, -7835, 2266, 7905, -2023, -7968, 1779, 8021, -1539, -8068, 1300, 8105, -1065, -8136, 831, 8159, -602, -8177, 374, 8186, -152, -8191, -69, 8189, 284, -8182, -497, 8168, 704, -8152, -909, 8128, 1108, -8102, -1304, 8070, 1494, -8036, -1681, 7996, 1862, -7955, -2041, 7909, 2212, -7863, -2382, 7811, 2544, -7760, -2704, 7704, 2857, -7648, -3008, 7589, 3152, -7531, -3293, 7469, 3428, -7408, -3561, 7345, 3687, -7283, -3811, 7219, 3928, -7156, -4043, 7092, 4152, -7029, -4258, 6965, 4359, -6904, -4457, 6841, 4550, -6781, -4640, 6720, 4725, -6662, -4808, 6602, 4885, -6547, -4961, 6490, 5031, -6437, -5099, 6384, 5162, -6335, -5224, 6285, 5280, -6239, -5335, 6193, 5385, -6151, -5434, 6109, 5477, -6071, -5520, 6034, 5558, -6000, -5594, 5967, 5626, -5939, -5657, 5911, 5683, -5887, -5708, 5864, 5729, -5845, -5749, 5827, 5764, -5813, -5778, 5800, 5788, -5792, -5797, 5784, 5801, -5781, -5805, 5778, 5804, -5780, -5803, 5783, 5797, -5790, -5790, 5798, 5779, -5811, -5767, 5824, 5750, -5842, -5733, 5860, 5711, -5883, -5688, 5906, 5660, -5934, -5632, 5962, 5599, -5995, -5564, 6028, 5525, -6065, -5485, 6103, 5440, -6144, -5394, 6186, 5343, -6232, -5290, 6277, 5232, -6327, -5173, 6376, 5109, -6429, -5043, 6482, 4971, -6538, -4898, 6593, 4820, -6652, -4739, 6710, 4653, -6771, -4565, 6831, 4471, -6894, -4376, 6955, 4274, -7019, -4170, 7082, 4060, -7146, -3947, 7209, 3829, -7273, -3708, 7335, 3580, -7398, -3451, 7459, 3314, -7521, -3176, 7580, 3030, -7639, -2882, 7695, 2728, -7751, -2571, 7803, 2407, -7855, -2241, 7902, 2068, -7948, -1892, 7990, 1710, -8030, -1525, 8065, 1334, -8097, -1140, 8124, 940, -8148, -738, 8166, 530, -8180, -319, 8188, 103, -8191, 115, 8187, -339, -8179, 565, 8162, -795, -8141, 1027, 8110, -1263, -8074, 1500, 8029, -1742, -7977, 1983, 7915, -2228, -7847, 2473, 7768, -2721, -7682, 2967, 7585, -3216, -7480, 3462, 7364, -3711, -7239, 3956, 7103, -4202, -6958, 4444, 6800, -4686, -6635, 4922, 6456, -5158, -6269, 5387, 6068, -5614, -5859, 5833, 5637, -6049, -5406, 6257, 5162, -6459, -4910, 6652, 4645, -6839, -4371, 7014, 4085, -7182, -3791, 7337, 3486, -7484, -3173, 7617, 2848, -7739, -2518, 7847, 2177, -7943, -1830, 8022, 1474, -8089, -1113, 8138, 745, -8172, -373, 8188, -5, -8189, 385, 8170, -770, -8135, 1155, 8079, -1542, -8006, 1928, 7911, -2315, -7798, 2698, 7664, -3080, -7511, 3456, 7336, -3828, -7142, 4191, 6926, -4549, -6692, 4896, 6436, -5234, -6161, 5559, 5865, -5873, -5551, 6170, 5217, -6454, -4867, 6719, 4496, -6968, -4112, 7196, 3709, -7405, -3293, 7590, 2862, -7754, -2419, 7892, 1963, -8006, -1499, 8093, 1024, -8154, -544, 8185, 57, -8189, 433, 8162, -927, -8107, 1419, 8019, -1911, -7903, 2398, 7753, -2881, -7575, 3354, 7363, -3820, -7122, 4271, 6848, -4710, -6547, 5131, 6214, -5536, -5854, 5917, 5465, -6278, -5052, 6612, 4611, -6920, -4149, 7198, 3663, -7447, -3158, 7661, 2634, -7842, -2096, 7986, 1542, -8094, -979, 8161, 406, -8191, 171, 8177, -753, -8125, 1333, 8028, -1911, -7891, 2482, 7710, -3044, -7489, 3592, 7223, -4126, -6919, 4638, 6573, -5130, -6190, 5594, 5767, -6031, -5311, 6433, 4819, -6803, -4299, 7133, 3747, -7424, -3172, 7669, 2572, -7872, -1955, 8025, 1320, -8130, -676, 8183, 21, -8186, 636, 8133, -1294, -8030, 1945, 7870, -2589, -7659, 3217, 7393, -3829, -7077, 4416, 6708, -4977, -6292, 5504, 5828, -5997, -5321, 6448, 4771, -6856, -4186, 7214, 3564, -7522, -2915, 7774, 2238, -7970, -1543, 8104, 830, -8178, -109, 8187, -618, -8133, 1342, 8011, -2061, -7827, 2766, 7576, -3453, -7264, 4113, 6888, -4743, -6454, 5336, 5961, -5887, -5417, 6389, 4822, -6840, -4183, 7231, 3503, -7561, -2790, 7824, 2047, -8020, -1284, 8141, 503, -8191, 284, 8162, -1074, -8059, 1856, 7877, -2626, -7622, 3372, 7289, -4091, -6886, 4771, 6412, -5409, -5874, 5995, 5273, -6525, -4619, 6989, 3912, -7386, -3164, 7706, 2377, -7950, -1565, 8109, 730, -8186, 114, 8173, -963, -8074, 1802, 7884, -2628, -7610, 3427, 7248, -4193, -6806, 4913, 6283, -5582, -5689, 6189, 5025, -6730, -4302, 7192, 3524, -7575, -2703, 7867, 1845, -8070, -964, 8174, 65, -8182, 836, 8089, -1733, -7898, 2610, 7606, -3460, -7220, 4268, 6739, -5028, -6173, 5724, 5524, -6352, -4803, 6898, 4015, -7358, -3173, 7721, 2283, -7985, -1362, 8142, 417, -8191, 535, 8128, -1486, -7955, 2418, 7669, -3323, -7278, 4182, 6782, -4988, -6190, 5724, 5506, -6383, -4742, 6951, 3905, -7423, -3010, 7786, 2066, -8037, -1089, 8169, 91, -8181, 910, 8068, -1904, -7835, 2869, 7479, -3797, -7009, 4667, 6426, -5470, -5743, 6188, 4966, -6814, -4109, 7331, 3181, -7735, -2201, 8013, 1180, -8165, -139, 8181, -911, -8065, 1948, 7813, -2957, -7432, 3919, 6922, -4820, -6295, 5640, 5557, -6369, -4723, 6988, 3803, -7490, -2815, 7861, 1772, -8097, -697, 8189, -397, -8137, 1485, 7937, -2552, -7595, 3574, 7111, -4537, -6497, 5417, 5760, -6202, -4916, 6873, 3974, -7418, -2957, 7824, 1879, -8084, -763, 8188, -373, -8137, 1504, 7927, -2610, -7563, 3668, 7048, -4659, -6393, 5558, 5608, -6352, -4710, 7019, 3712, -7548, -2638, 7923, 1505, -8139, -339, 8187, -840, -8067, 2002, 7776, -3129, -7324, 4191, 6713, -5170, -5960, 6039, 5075, -6784, -4081, 7383, 2993, -7825, -1838, 8096, 638, -8191, 578, 8104, -1787, -7839, 2957, 7395, -4067, -6785, 5086, 6018, -5995, -5113, 6768, 4087, -7389, -2965, 7839, 1769, -8110, -530, 8190, -727, -8079, 1968, 7775, -3168, -7287, 4295, 6620, -5323, -5794, 6223, 4823, -6977, -3734, 7560, 2548, -7961, -1298, 8164, 10, -8167, 1280, 7963, -2544, -7560, 3744, 6963, -4856, -6188, 5844, 5252, -6687, -4179, 7358, 2993, -7842, -1728, 8120, 412, -8188, 917, 8037, -2227, -7675, 3479, 7105, -4643, -6345, 5684, 5409)    
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L15�33_i
    );

    L21_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-8189, -444, 8116, 1755, -7833, -3020, 7345, 4202, -6670, -5276, 5822, 6209, -4828, -6983, 3710, 7575, -2502, -7975, 1230, 8170, 68, -8160, -1364, 7943, 2621, -7529, -3812, 6926, 4904, -6154, -5874, 5230, 6695, -4180, -7351, 3027, 7824, -1805, -8107, 539, 8190, 735, -8076, -1991, 7766, 3195, -7272, -4321, 6603, 5340, -5780, -6232, 4820, 6973, -3749, -7549, 2591, 7945, -1376, -8157, 129, 8176, 1116, -8007, -2335, 7651, 3495, -7122, -4575, 6429, 5546, -5593, -6390, 4629, 7086, -3564, -7622, 2420, 7984, -1225, -8168, 4, 8168, 1213, -7988, -2403, 7630, 3535, -7107, -4588, 6427, 5538, -5610, -6366, 4671, 7053, -3635, -7588, 2521, 7957, -1356, -8156, 164, 8179, 1028, -8030, -2197, 7710, 3315, -7230, -4364, 6598, 5316, -5832, -6158, 4943, 6869, -3957, -7438, 2889, 7851, -1767, -8105, 608, 8190, 558, -8112, -1712, 7868, 2827, -7468, -3885, 6918, 4862, -6233, -5741, 5424, 6503, -4512, -7137, 3511, 7627, -2446, -7970, 1333, 8154, -199, -8183, -938, 8052, 2053, -7769, -3128, 7336, 4139, -6767, -5071, 6069, 5903, -5260, -6625, 4353, 7219, -3369, -7679, 2322, 7994, -1237, -8163, 129, 8179, 976, -8049, -2063, 7770, 3108, -7353, -4096, 6802, 5007, -6133, -5828, 5354, 6541, -4484, -7138, 3535, 7607, -2527, -7942, 1476, 8136, -403, -8190, -676, 8101, 1738, -7874, -2771, 7510, 3751, -7022, -4668, 6413, 5501, -5699, -6241, 4890, 6873, -4002, -7391, 3049, 7782, -2048, -8046, 1015, 8176, 30, -8173, -1075, 8035, 2097, -7769, -3085, 7376, 4019, -6869, -4889, 6251, 5676, -5537, -6373, 4735, 6967, -3863, -7451, 2930, 7816, -1957, -8061, 953, 8178, 60, -8172, -1072, 8038, 2064, -7785, -3023, 7412, 3932, -6931, -4782, 6345, 5557, -5668, -6248, 4907, 6844, -4077, -7339, 3188, 7723, -2256, -7996, 1292, 8151, -314, -8190, -668, 8109, 1636, -7914, -2580, 7606, 3484, -7194, -4337, 6679, 5126, -6075, -5843, 5386, 6476, -4627, -7020, 3803, 7464, -2933, -7807, 2022, 8041, -1089, -8168, 142, 8184, 803, -8092, -1737, 7891, 2642, -7589, -3513, 7186, 4334, -6692, -5097, 6111, 5791, -5455, -6410, 4729, 6944, -3946, -7390, 3113, 7739, -2246, -7991, 1350, 8141, -442, -8191, -470, 8138, 1372, -7987, -2257, 7737, 3110, -7395, -3925, 6963, 4688, -6450, -5394, 5860, 6033, -5204, -6600, 4486, 7085, -3720, -7489, 2910, 7802, -2071, -8025, 1209, 8154, -337, -8191, -538, 8133, 1403, -7985, -2251, 7745, 3069, -7422, -3853, 7015, 4590, -6534, -5276, 5981, 5900, -5367, -6460, 4693, 6947, -3974, -7359, 3212, 7690, -2420, -7940, 1603, 8104, -774, -8184, -63, 8176, 895, -8086, -1717, 7911, 2517, -7658, -3290, 7326, 4026, -6922, -4721, 6449, 5365, -5915, -5955, 5321, 6483, -4679, -6947, 3992, 7340, -3270, -7662, 2516, 7908, -1743, -8080, 954, 8172, -160, -8188, -635, 8126, 1419, -7990, -2190, 7778, 2936, -7498, -3654, 7148, 4335, -6736, -4976, 6263, 5568, -5737, -6111, 5160, 6596, -4541, -7023, 3883, 7385, -3195, -7684, 2479, 7913, -1747, -8075, 1000, 8167, -249, -8191, -504, 8143, 1247, -8031, -1980, 7850, 2692, -7607, -3381, 7300, 4038, -6938, -4663, 6519, 5245, -6051, -5786, 5535, 6277, -4978, -6719, 4383, 7105, -3758, -7437, 3104, 7708, -2431, -7921, 1739, 8072, -1039, -8163, 332, 8190, 373, -8159, -1075, 8066, 1765, -7916, -2441, 7708, 3095, -7446, -3726, 7130, 4327, -6767, -4896, 6356, 5427, -5903, -5920, 5410, 6369, -4883, -6774, 4322, 7129, -3736, -7437, 3126, 7692, -2499, -7896, 1856, 8046, -1205, -8145, 546, 8188, 111, -8180, -767, 8117, 1413, -8006, -2050, 7842, 2670, -7633, -3272, 7374, 3850, -7074, -4404, 6729, 4927, -6347, -5421, 5927, 5877, -5475, -6299, 4990, 6681, -4480, -7024, 3945, 7322, -3391, -7580, 2817, 7791, -2232, -7960, 1636, 8081, -1034, -8159, 427, 8190, 177, -8177, -780, 8119, 1374, -8020, -1960, 7876, 2532, -7694, -3089, 7470, 3626, -7210, -4144, 6912, 4637, -6583, -5106, 6220, 5545, -5830, -5957, 5410, 6335, -4968, -6683, 4501, 6995, -4017, -7274, 3514, 7515, -2998, -7721, 2469, 7889, -1933, -8021, 1389, 8114, -842, -8172, 293, 8190, 254, -8175, -798, 8121, 1335, -8033, -1865, 7910, 2383, -7755, -2890, 7566, 3380, -7348, -3856, 7099, 4311, -6823, -4749, 6519, 5163, -6192, -5556, 5840, 5923, -5469, -6267, 5076, 6583, -4667, -6874, 4240, 7135, -3801, -7369, 3349, 7573, -2888, -7750, 2417, 7895, -1941, -8013, 1459, 8099, -976, -8159, 491, 8187, -8, -8188, -474, 8159, 950, -8105, -1423, 8022, 1886, -7914, -2342, 7779, 2786, -7621, -3220, 7437, 3640, -7233, -4048, 7005, 4438, -6758, -4815, 6490, 5173, -6206, -5516, 5902, 5837, -5585, -6142, 5251, 6425, -4906, -6689, 4547, 6931, -4179, -7154, 3799, 7354, -3413, -7534, 3018, 7690, -2619, -7827, 2214, 7940, -1807, -8033, 1396, 8103, -986, -8154, 574, 8182, -165, -8191, -244, 8178, 648, -8147, -1049, 8095, 1443, -8026, -1834, 7936, 2215, -7831, -2591, 7706, 2957, -7567, -3315, 7410, 3662, -7239, -4001, 7053, 4326, -6854, -4643, 6640, 4945, -6416, -5237, 6178, 5514, -5932, -5781, 5673, 6032, -5407, -6271, 5131, 6495, -4848, -6707, 4557, 6902, -4261, -7086, 3958, 7253, -3651, -7408, 3339, 7547, -3025, -7674, 2706, 7784, -2387, -7883, 2065, 7966, -1743, -8037, 1420, 8093, -1098, -8138, 776, 8167, -456, -8186, 137, 8190, 178, -8185, -492, 8165, 801, -8136, -1108, 8093, 1409, -8042, -1708, 7978, 1999, -7906, -2288, 7822, 2569, -7731, -2846, 7629, 3115, -7520, -3380, 7401, 3637, -7276, -3888, 7141, 4131, -7002, -4369, 6854, 4598, -6701, -4822, 6541, 5036, -6377, -5245, 6206, 5444, -6032, -5638, 5852, 5822, -5670, -6000, 5482, 6169, -5293, -6333, 5098, 6486, -4903, -6635, 4704, 6774, -4505, -6907, 4302, 7031, -4099, -7150, 3893, 7260, -3689, -7365, 3482, 7461, -3276, -7552, 3068, 7635, -2863, -7713, 2655, 7782, -2451, -7848, 2245, 7905, -2042, -7958, 1838, 8004, -1638, -8046, 1437, 8080, -1240, -8112, 1043, 8136, -849, -8157, 656, 8171, -467, -8183, 278, 8188, -94, -8191, -90, 8189, 269, -8184, -448, 8173, 622, -8161, -794, 8143, 962, -8124, -1129, 8101, 1291, -8076, -1452, 8046, 1608, -8016, -1762, 7982, 1912, -7947, -2060, 7908, 2203, -7869, -2345, 7827, 2481, -7785, -2617, 7739, 2747, -7694, -2876, 7645, 3000, -7598, -3122, 7547, 3240, -7498, -3356, 7446, 3467, -7395, -3577, 7342, 3682, -7291, -3786, 7237, 3885, -7185, -3983, 7131, 4076, -7079, -4167, 7025, 4255, -6973, -4341, 6920, 4422, -6869, -4503, 6817, 4578, -6767, -4654, 6716, 4724, -6667, -4794, 6617, 4859, -6570, -4924, 6523, 4984, -6478, -5043, 6432, 5099, -6389, -5154, 6345, 5204, -6305, -5254, 6264, 5300, -6226, -5346, 6188, 5387, -6153, -5428, 6117, 5465, -6085, -5502, 6052, 5535, -6023, -5568, 5994, 5596, -5968, -5625, 5942, 5650, -5919, -5674, 5896, 5695, -5877, -5716, 5858, 5733, -5842, -5750, 5826, 5763, -5814, -5776, 5802, 5786, -5794, -5795, 5785, 5801, -5780, -5807, 5775, 5809, -5774, -5811, 5772, 5810, -5775, -5808, 5777, 5803, -5783, -5798, 5789, 5789, -5799, -5781, 5809, 5768, -5822, -5756, 5835, 5739, -5852, -5723, 5869, 5703, -5890, -5683, 5910, 5659, -5934, -5635, 5957, 5607, -5984, -5579, 6011, 5547, -6042, -5515, 6072, 5479, -6105, -5443, 6138, 5402, -6175, -5362, 6211, 5317, -6250, -5272, 6289, 5223, -6331, -5173, 6372, 5119, -6416, -5065, 6459, 5006, -6506, -4947, 6552, 4883, -6600, -4819, 6647, 4750, -6698, -4681, 6747, 4607, -6798, -4532, 6849, 4453, -6901, -4372, 6952, 4287, -7006, -4201, 7058, 4110, -7112, -4019, 7164, 3922, -7218, -3824, 7270, 3721, -7323, -3618, 7375, 3509, -7428, -3399, 7478, 3284, -7529, -3168, 7578, 3046, -7628, -2924, 7675, 2796, -7723, -2667, 7767, 2533, -7812, -2397, 7853, 2257, -7894, -2115, 7932, 1968, -7969, -1820, 8003, 1666, -8036, -1512, 8064, 1352, -8092, -1191, 8115, 1026, -8137, -859, 8154, 687, -8169, -514, 8179, 337, -8188, -159, 8190, -24, -8191, 207, 8185, -395, -8177, 583, 8162, -776, -8145, 969, 8121, -1165, -8093, 1362, 8059, -1562, -8021, 1762, 7976, -1965, -7927, 2168, 7870, -2373, -7809, 2578, 7739, -2785, -7666, 2990, 7584, -3198, -7497, 3403, 7402, -3611, -7302, 3816, 7192, -4022, -7078, 4225, 6955, -4428, -6826, 4628, 6688, -4829, -6544, 5024, 6391, -5220, -6233, 5410, 6065, -5599, -5891, 5783, 5708, -5965, -5519, 6140, 5320, -6313, -5116, 6479, 4903, -6642, -4684, 6796, 4456, -6947, -4223, 7089, 3981, -7226, -3733, 7354, 3478, -7476, -3217, 7588, 2948, -7694, -2675, 7788, 2394, -7876, -2110, 7951, 1818, -8019, -1523, 8075, 1222, -8121, -918, 8155, 609, -8179, -298, 8189, -18, -8190, 334, 8176, -655, -8151, 975, 8111, -1298, -8060, 1620, 7994, -1944, -7917, 2265, 7823, -2586, -7718, 2904, 7596, -3221, -7463, 3533, 7313, -3843, -7151, 4146, 6973, -4446, -6783, 4738, 6576, -5025, -6358, 5303, 6124, -5574, -5878, 5834, 5616, -6087, -5344, 6327, 5057, -6557, -4759, 6774, 4447, -6979, -4126, 7170, 3791, -7348, -3448, 7509, 3093, -7656, -2731, 7785, 2358, -7899, -1979, 7993, 1592, -8072, -1199, 8129, 800, -8170, -398, 8188, -10, -8189, 418, 8167, -830, -8126, 1240, 8062, -1652, -7978, 2060, 7872, -2466, -7745, 2867, 7595, -3265, -7425, 3653, 7232, -4036, -7019, 4408, 6783, -4772, -6528, 5122, 6251, -5461, -5956, 5784, 5639, -6093, -5306, 6384, 4952, -6659, -4584, 6913, 4197, -7149, -3797, 7362, 3380, -7554, -2952, 7721, 2510, -7866, -2060, 7983, 1598, -8077, -1131, 8142, 655, -8181, -176, 8190, -308, -8173, 792, 8125, -1277, -8050, 1758, 7943, -2238, -7809, 2710, 7643, -3176, -7450, 3631, 7227, -4076, -6976, 4506, 6696, -4923, -6390, 5321, 6056, -5702, -5699, 6061, 5314, -6399, -4909, 6710, 4479, -6998, -4031, 7256, 3562, -7488, -3078, 7687, 2576, -7856, -2063, 7990, 1536, -8092, -1003, 8158, 460, -8189, 85, 8183, -634, -8141, 1182, 8060, -1728, -7944, 2267, 7789, -2800, -7598, 3320, 7369, -3829, -7105, 4319, 6804, -4794, -6471, 5245, 6103, -5674, -5705, 6075, 5275, -6450, -4818, 6791, 4333, -7102, -3826, 7375, 3294, -7614, -2745, 7811, 2178, -7971, -1598, 8086, 1005, -8161, -407, 8190, -199, -8176, 804, 8115, -1409, -8011, 2007, 7860, -2598, -7666, 3175, 7425, -3738, -7142, 4279, 6815, -4801, -6449, 5294, 6041, -5760, -5598, 6191, 5118, -6589, -4606, 6947, 4063, -7266, -3495, 7539, 2900, -7769, -2287, 7949, 1656, -8082, -1013, 8162, 360, -8191, 297, 8166, -956, -8090, 1610, 7959, -2257, -7776, 2890, 7539, -3508, -7252, 4103, 6914, -4674, -6528, 5213, 6095, -5721, -5619, 6189, 5101, -6617, -4547, 6998, 3957, -7333, -3338, 7615, 2691, -7844, -2024, 8016, 1337, -8131, -641, 8185, -65, -8181, 771, 8113, -1476, -7986, 2170, 7795, -2852, -7547, 3513, 7237, -4151, -6872, 4756, 6451, -5329, -5978, 5860, 5455, -6348, -4889, 6785, 4279, -7170, -3634, 7497, 2956, -7766, -2252, 7969, 1526, -8109, -787, 8180, 36, -8184, 715, 8118, -1465, -7983, 2203, 7778, -2927, -7506, 3625, 7167, -4296, -6765, 4930, 6301, -5525, -5781, 6070, 5206, -6564, -4584, 6999, 3916, -7373, -3212, 7680, 2475, -7918, -1714, 8083, 933, -8174, -142, 8187, -654, -8124, 1445, 7982, -2226, -7765, 2987, 7470, -3723, -7104, 4423, 6666, -5084, -6163, 5696, 5595, -6254, -4972, 6750, 4294, -7182, -3574, 7540, 2813, -7825, -2023, 8029, 1208, -8153, -380, 8190, -457, -8145, 1290, 8011, -2113, -7795, 2915, 7493, -3690, -7113, 4426, 6652, -5118, -6121, 5755, 5519, -6333, -4857, 6841, 4137, -7278, -3371, 7632, 2564, -7905, -1727, 8087, 867, -8180, 4, 8179, -880, -8085, 1746, 7897, -2596, -7618, 3417, 7248, -4202, -6794, 4938, 6256, -5620, -5645, 6235, 4962, -6779, -4221, 7241, 3424, -7619, -2585, 7903, 1710, -8093, -814, 8183, -97, -8173, 1007, 8059, -1909, -7847, 2788, 7532, -3636, -7124, 4438, 6622, -5188, -6036, 5871, 5368, -6482, -4631, 7009, 3830, -7448, -2978, 7788, 2083, -8029, -1160, 8161, 216, -8187, 730, 8102, -1672, -7908, 2591, 7605, -3479, -7200, 4321, 6693, -5107, -6094, 5823, 5407, -6462, -4645, 7010, 3813, -7463, -2928, 7810, 1997, -8049, -1037, 8172, 58, -8180, 922, 8068, -1894, -7841, 2839, 7497, -3747, -7044, 4600, 6485, -5389, -5830, 6099, 5084, -6721, -4263, 7242, 3373, -7658, -2433, 7956, 1450, -8136, -446, 8190, -571, -8120, 1579, 7923, -2567, -7604, 3515, 7163, -4413, -6611, 5242, 5951, -5992, -5197, 6646, 4357, -7198, -3447, 7634, 2476, -7950, -1466, 8135, 427, -8191, 619, 8111, -1660, -7898, 2674, 7553, -3648, -7084, 4562, 6493, -5403, -5793, 6154, 4993, -6805, -4108, 7339, 3148, -7752, -2135, 8030, 1080, -8173, -7, 8173, -1072, -8033, 2132, 7749, -3160, -7332, 4132, 6781, -5035, -6111, 5850, 5329, -6563, -4452, 7159, 3490, -7628, -2465, 7959, 1391, -8148, -291, 8186, -819, -8076, 1914, 7815, -2979, -7410, 3988, 6865, -4928, -6191, 5775, 5398, -6517, -4503, 7136, 3519, -7622, -2467, 7962, 1363, -8152, -233, 8184, -906, -8059, 2028, 7774, -3115, -7340, 4141, 6758, -5091, -6044, 5940, 5207, -6675, -4266, 7276, 3236, -7735, -2140, 8038, 998, -8181, 166, 8156, -1331, -7967, 2469, 7612, -3561, -7103, 4580, 6443, -5509, -5650, 6323, 4736, -7008, -3723, 7547, 2627, -7929, -1475, 8143, 288, -8186, 906, 8052, -2085, -7748, 3220, 7274, -4290, -6644, 5267, 5867, -6134, -4962, 6866, 3944, -7452, -2840, 7872, 1668, -8122, -459, 8189, -764, -8076, 1972, 7779, -3139, -7309, 4236, 6671, -5242, -5882, 6128, 4956, -6878, -3916, 7470, 2782, -7894, -1583, 8133, 343, -8187, 905, 8047, -2136, -7721, 3319, 7211, -4427, -6532, 5431, 5694, -6310, -4721, 7038, 3632, -7601, -2455, 7981, 1215, -8171, 56, 8161, -1329, -7955, 2571, 7552, -3754, -6964, 4845, 6203, -5821, -5288, 6653, 4238, -7322, -3083, 7809, 1846, -8102, -562, 8190, -741, -8073, 2025, 7749, -3262, -7230, 4417, 6522, -5462, -5647, 6367, 4623, -7112, -3480, 7671, 2242, -8034, -945, 8186, -382, -8125, 1699, 7848, -2975, -7365, 4173, 6684, -5265, -5825, 6216, 4807, -7004, -3660, 7603, 2410, -8001, -1094)    
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L21_i
    );

    L21C31_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (8188, 443, -8117, -1756, 7832, 3019, -7346, -4203, 6669, 5275, -5823, -6210, 4827, 6982, -3711, -7576, 2501, 7974, -1231, -8171, -69, 8159, 1363, -7944, -2622, 7528, 3811, -6927, -4905, 6153, 5873, -5231, -6696, 4179, 7350, -3028, -7825, 1804, 8106, -540, -8191, -736, 8075, 1990, -7767, -3196, 7271, 4320, -6604, -5341, 5779, 6231, -4821, -6974, 3748, 7548, -2592, -7946, 1375, 8156, -130, -8177, -1117, 8006, 2334, -7652, -3496, 7121, 4574, -6430, -5547, 5592, 6389, -4630, -7087, 3563, 7621, -2421, -7985, 1224, 8167, -5, -8169, -1214, 7987, 2402, -7631, -3536, 7106, 4587, -6428, -5539, 5609, 6365, -4672, -7054, 3634, 7587, -2522, -7958, 1355, 8155, -165, -8180, -1029, 8029, 2196, -7711, -3316, 7229, 4363, -6599, -5317, 5831, 6157, -4944, -6870, 3956, 7437, -2890, -7852, 1766, 8104, -609, -8191, -559, 8111, 1711, -7869, -2828, 7467, 3884, -6919, -4863, 6232, 5740, -5425, -6504, 4511, 7136, -3512, -7628, 2445, 7969, -1334, -8155, 198, 8182, 937, -8053, -2054, 7768, 3127, -7337, -4140, 6766, 5070, -6070, -5904, 5259, 6624, -4354, -7220, 3368, 7678, -2323, -7995, 1236, 8162, -130, -8180, -977, 8048, 2062, -7771, -3109, 7352, 4095, -6803, -5008, 6132, 5827, -5355, -6542, 4483, 7137, -3536, -7608, 2526, 7941, -1477, -8137, 402, 8189, 675, -8102, -1739, 7873, 2770, -7511, -3752, 7021, 4667, -6414, -5502, 5698, 6240, -4891, -6874, 4001, 7390, -3050, -7783, 2047, 8045, -1016, -8177, -31, 8172, 1074, -8036, -2098, 7768, 3084, -7377, -4020, 6868, 4888, -6252, -5677, 5536, 6372, -4736, -6968, 3862, 7450, -2931, -7817, 1956, 8060, -954, -8179, -61, 8171, 1071, -8039, -2065, 7784, 3022, -7413, -3933, 6930, 4781, -6346, -5558, 5667, 6247, -4908, -6845, 4076, 7338, -3189, -7724, 2255, 7995, -1293, -8152, 313, 8189, 667, -8110, -1637, 7913, 2579, -7607, -3485, 7193, 4336, -6680, -5127, 6074, 5842, -5387, -6477, 4626, 7019, -3804, -7465, 2932, 7806, -2023, -8042, 1088, 8167, -143, -8185, -804, 8091, 1736, -7892, -2643, 7588, 3512, -7187, -4335, 6691, 5096, -6112, -5792, 5454, 6409, -4730, -6945, 3945, 7389, -3114, -7740, 2245, 7990, -1351, -8142, 441, 8190, 469, -8139, -1373, 7986, 2256, -7738, -3111, 7394, 3924, -6964, -4689, 6449, 5393, -5861, -6034, 5203, 6599, -4487, -7086, 3719, 7488, -2911, -7803, 2070, 8024, -1210, -8155, 336, 8190, 537, -8134, -1404, 7984, 2250, -7746, -3070, 7421, 3852, -7016, -4591, 6533, 5275, -5982, -5901, 5366, 6459, -4694, -6948, 3973, 7358, -3213, -7691, 2419, 7939, -1604, -8105, 773, 8183, 62, -8177, -896, 8085, 1716, -7912, -2518, 7657, 3289, -7327, -4027, 6921, 4720, -6450, -5366, 5914, 5954, -5322, -6484, 4678, 6946, -3993, -7341, 3269, 7661, -2517, -7909, 1742, 8079, -955, -8173, 159, 8187, 634, -8127, -1420, 7989, 2189, -7779, -2937, 7497, 3653, -7149, -4336, 6735, 4975, -6264, -5569, 5736, 6110, -5161, -6597, 4540, 7022, -3884, -7386, 3194, 7683, -2480, -7914, 1746, 8074, -1001, -8168, 248, 8190, 503, -8144, -1248, 8030, 1979, -7851, -2693, 7606, 3380, -7301, -4039, 6937, 4662, -6520, -5246, 6050, 5785, -5536, -6278, 4977, 6718, -4384, -7106, 3757, 7436, -3105, -7709, 2430, 7920, -1740, -8073, 1038, 8162, -333, -8191, -374, 8158, 1074, -8067, -1766, 7915, 2440, -7709, -3096, 7445, 3725, -7131, -4328, 6766, 4895, -6357, -5428, 5902, 5919, -5411, -6370, 4882, 6773, -4323, -7130, 3735, 7436, -3127, -7693, 2498, 7895, -1857, -8047, 1204, 8144, -547, -8189, -112, 8179, 766, -8118, -1414, 8005, 2049, -7843, -2671, 7632, 3271, -7375, -3851, 7073, 4403, -6730, -4928, 6346, 5420, -5928, -5878, 5474, 6298, -4991, -6682, 4479, 7023, -3946, -7323, 3390, 7579, -2818, -7792, 2231, 7959, -1637, -8082, 1033, 8158, -428, -8191, -178, 8176, 779, -8120, -1375, 8019, 1959, -7877, -2533, 7693, 3088, -7471, -3627, 7209, 4143, -6913, -4638, 6582, 5105, -6221, -5546, 5829, 5956, -5411, -6336, 4967, 6682, -4502, -6996, 4016, 7273, -3515, -7516, 2997, 7720, -2470, -7890, 1932, 8020, -1390, -8115, 841, 8171, -294, -8191, -255, 8174, 797, -8122, -1336, 8032, 1864, -7911, -2384, 7754, 2889, -7567, -3381, 7347, 3855, -7100, -4312, 6822, 4748, -6520, -5164, 6191, 5555, -5841, -5924, 5468, 6266, -5077, -6584, 4666, 6873, -4241, -7136, 3800, 7368, -3350, -7574, 2887, 7749, -2418, -7896, 1940, 8012, -1460, -8100, 975, 8158, -492, -8188, 7, 8187, 473, -8160, -951, 8104, 1422, -8023, -1887, 7913, 2341, -7780, -2787, 7620, 3219, -7438, -3641, 7232, 4047, -7006, -4439, 6757, 4814, -6491, -5174, 6205, 5515, -5903, -5838, 5584, 6141, -5252, -6426, 4905, 6688, -4548, -6932, 4178, 7153, -3800, -7355, 3412, 7533, -3019, -7691, 2618, 7826, -2215, -7941, 1806, 8032, -1397, -8104, 985, 8153, -575, -8183, 164, 8190, 243, -8179, -649, 8146, 1048, -8096, -1444, 8025, 1833, -7937, -2216, 7830, 2590, -7707, -2958, 7566, 3314, -7411, -3663, 7238, 4000, -7054, -4327, 6853, 4642, -6641, -4946, 6415, 5236, -6179, -5515, 5931, 5780, -5674, -6033, 5406, 6270, -5132, -6496, 4847, 6706, -4558, -6903, 4260, 7085, -3959, -7254, 3650, 7407, -3340, -7548, 3024, 7673, -2707, -7785, 2386, 7882, -2066, -7967, 1742, 8036, -1421, -8094, 1097, 8137, -777, -8168, 455, 8185, -138, -8191, -179, 8184, 491, -8166, -802, 8135, 1107, -8094, -1410, 8041, 1707, -7979, -2000, 7905, 2287, -7823, -2570, 7730, 2845, -7630, -3116, 7519, 3379, -7402, -3638, 7275, 3887, -7142, -4132, 7001, 4368, -6855, -4599, 6700, 4821, -6542, -5037, 6376, 5244, -6207, -5445, 6031, 5637, -5853, -5823, 5669, 5999, -5483, -6170, 5292, 6332, -5099, -6487, 4902, 6634, -4705, -6775, 4504, 6906, -4303, -7032, 4098, 7149, -3894, -7261, 3688, 7364, -3483, -7462, 3275, 7551, -3069, -7636, 2862, 7712, -2656, -7783, 2450, 7847, -2246, -7906, 2041, 7957, -1839, -8005, 1637, 8045, -1438, -8081, 1239, 8111, -1044, -8137, 848, 8156, -657, -8172, 466, 8182, -279, -8189, 93, 8190, 89, -8190, -270, 8183, 447, -8174, -623, 8160, 793, -8144, -963, 8123, 1128, -8102, -1292, 8075, 1451, -8047, -1609, 8015, 1761, -7983, -1913, 7946, 2059, -7909, -2204, 7868, 2344, -7828, -2482, 7784, 2616, -7740, -2748, 7693, 2875, -7646, -3001, 7597, 3121, -7548, -3241, 7497, 3355, -7447, -3468, 7394, 3576, -7343, -3683, 7290, 3785, -7238, -3886, 7184, 3982, -7132, -4077, 7078, 4166, -7026, -4256, 6972, 4340, -6921, -4423, 6868, 4502, -6818, -4579, 6766, 4653, -6717, -4725, 6666, 4793, -6618, -4860, 6569, 4923, -6524, -4985, 6477, 5042, -6433, -5100, 6388, 5153, -6346, -5205, 6304, 5253, -6265, -5301, 6225, 5345, -6189, -5388, 6152, 5427, -6118, -5466, 6084, 5501, -6053, -5536, 6022, 5567, -5995, -5597, 5967, 5624, -5943, -5651, 5918, 5673, -5897, -5696, 5876, 5715, -5859, -5734, 5841, 5749, -5827, -5764, 5813, 5775, -5803, -5787, 5793, 5794, -5786, -5802, 5779, 5806, -5776, -5810, 5773, 5810, -5773, -5811, 5774, 5807, -5778, -5804, 5782, 5797, -5790, -5790, 5798, 5780, -5810, -5769, 5821, 5755, -5836, -5740, 5851, 5722, -5870, -5704, 5889, 5682, -5911, -5660, 5933, 5634, -5958, -5608, 5983, 5578, -6012, -5548, 6041, 5514, -6073, -5480, 6104, 5442, -6139, -5403, 6174, 5361, -6212, -5318, 6249, 5271, -6290, -5224, 6330, 5172, -6373, -5120, 6415, 5064, -6460, -5007, 6505, 4946, -6553, -4884, 6599, 4818, -6648, -4751, 6697, 4680, -6748, -4608, 6797, 4531, -6850, -4454, 6900, 4371, -6953, -4288, 7005, 4200, -7059, -4111, 7111, 4018, -7165, -3923, 7217, 3823, -7271, -3722, 7322, 3617, -7376, -3510, 7427, 3398, -7479, -3285, 7528, 3167, -7579, -3047, 7627, 2923, -7676, -2797, 7722, 2666, -7768, -2534, 7811, 2396, -7854, -2258, 7893, 2114, -7933, -1969, 7968, 1819, -8004, -1667, 8035, 1511, -8065, -1353, 8091, 1190, -8116, -1027, 8136, 858, -8155, -688, 8168, 513, -8180, -338, 8187, 158, -8191, 23, 8190, -208, -8186, 394, 8176, -584, -8163, 775, 8144, -970, -8122, 1164, 8092, -1363, -8060, 1561, 8020, -1763, -7977, 1964, 7926, -2169, -7871, 2372, 7808, -2579, -7740, 2784, 7665, -2991, -7585, 3197, 7496, -3404, -7403, 3610, 7301, -3817, -7193, 4021, 7077, -4226, -6956, 4427, 6825, -4629, -6689, 4828, 6543, -5025, -6392, 5219, 6232, -5411, -6066, 5598, 5890, -5784, -5709, 5964, 5518, -6141, -5321, 6312, 5115, -6480, -4904, 6641, 4683, -6797, -4457, 6946, 4222, -7090, -3982, 7225, 3732, -7355, -3479, 7475, 3216, -7589, -2949, 7693, 2674, -7789, -2395, 7875, 2109, -7952, -1819, 8018, 1522, -8076, -1223, 8120, 917, -8156, -610, 8178, 297, -8190, 17, 8189, -335, -8177, 654, 8150, -976, -8112, 1297, 8059, -1621, -7995, 1943, 7916, -2266, -7824, 2585, 7717, -2905, -7597, 3220, 7462, -3534, -7314, 3842, 7150, -4147, -6974, 4445, 6782, -4739, -6577, 5024, 6357, -5304, -6125, 5573, 5877, -5835, -5617, 6086, 5343, -6328, -5058, 6556, 4758, -6775, -4448, 6978, 4125, -7171, -3792, 7347, 3447, -7510, -3094, 7655, 2730, -7786, -2359, 7898, 1978, -7994, -1593, 8071, 1198, -8130, -801, 8169, 397, -8189, 9, 8188, -419, -8168, 829, 8125, -1241, -8063, 1651, 7977, -2061, -7873, 2465, 7744, -2868, -7596, 3264, 7424, -3654, -7233, 4035, 7018, -4409, -6784, 4771, 6527, -5123, -6252, 5460, 5955, -5785, -5640, 6092, 5305, -6385, -4953, 6658, 4583, -6914, -4198, 7148, 3796, -7363, -3381, 7553, 2951, -7722, -2511, 7865, 2059, -7984, -1599, 8076, 1130, -8143, -656, 8180, 175, -8191, 307, 8172, -793, -8126, 1276, 8049, -1759, -7944, 2237, 7808, -2711, -7644, 3175, 7449, -3632, -7228, 4075, 6975, -4507, -6697, 4922, 6389, -5322, -6057, 5701, 5698, -6062, -5315, 6398, 4908, -6711, -4480, 6997, 4030, -7257, -3563, 7487, 3077, -7688, -2577, 7855, 2062, -7991, -1537, 8091, 1002, -8159, -461, 8188, -86, -8184, 633, 8140, -1183, -8061, 1727, 7943, -2268, -7790, 2799, 7597, -3321, -7370, 3828, 7104, -4320, -6805, 4793, 6470, -5246, -6104, 5673, 5704, -6076, -5276, 6449, 4817, -6792, -4334, 7101, 3825, -7376, -3295, 7613, 2744, -7812, -2179, 7970, 1597, -8087, -1006, 8160, 406, -8191, 198, 8175, -805, -8116, 1408, 8010, -2008, -7861, 2597, 7665, -3176, -7426, 3737, 7141, -4280, -6816, 4800, 6448, -5295, -6042, 5759, 5597, -6192, -5119, 6588, 4605, -6948, -4064, 7265, 3494, -7540, -2901, 7768, 2286, -7950, -1657, 8081, 1012, -8163, -361, 8190, -298, -8167, 955, 8089, -1611, -7960, 2256, 7775, -2891, -7540, 3507, 7251, -4104, -6915, 4673, 6527, -5214, -6096, 5720, 5618, -6190, -5102, 6616, 4546, -6999, -3958, 7332, 3337, -7616, -2692, 7843, 2023, -8017, -1338, 8130, 640, -8186, 64, 8180, -772, -8114, 1475, 7985, -2171, -7796, 2851, 7546, -3514, -7238, 4150, 6871, -4757, -6452, 5328, 5977, -5861, -5456, 6347, 4888, -6786, -4280, 7169, 3633, -7498, -2957, 7765, 2251, -7970, -1527, 8108, 786, -8181, -37, 8183, -716, -8119, 1464, 7982, -2204, -7779, 2926, 7505, -3626, -7168, 4295, 6764, -4931, -6302, 5524, 5780, -6071, -5207, 6563, 4583, -7000, -3917, 7372, 3211, -7681, -2476, 7917, 1713, -8084, -934, 8173, 141, -8188, 653, 8123, -1446, -7983, 2225, 7764, -2988, -7471, 3722, 7103, -4424, -6667, 5083, 6162, -5697, -5596, 6253, 4971, -6751, -4295, 7181, 3573, -7541, -2814, 7824, 2022, -8030, -1209, 8152, 379, -8191, 456, 8144, -1291, -8012, 2112, 7794, -2916, -7494, 3689, 7112, -4427, -6653, 5117, 6120, -5756, -5520, 6332, 4856, -6842, -4138, 7277, 3370, -7633, -2565, 7904, 1726, -8088, -868, 8179, -5, -8180, 879, 8084, -1747, -7898, 2595, 7617, -3418, -7249, 4201, 6793, -4939, -6257, 5619, 5644, -6236, -4963, 6778, 4220, -7242, -3425, 7618, 2584, -7904, -1711, 8092, 813, -8184, 96, 8172, -1008, -8060, 1908, 7846, -2789, -7533, 3635, 7123, -4439, -6623, 5187, 6035, -5872, -5369, 6481, 4630, -7010, -3831, 7447, 2977, -7789, -2084, 8028, 1159, -8162, -217, 8186, -731, -8103, 1671, 7907, -2592, -7606, 3478, 7199, -4322, -6694, 5106, 6093, -5824, -5408, 6461, 4644, -7011, -3814, 7462, 2927, -7811, -1998, 8048, 1036, -8173, -59, 8179, -923, -8069, 1893, 7840, -2840, -7498, 3746, 7043, -4601, -6486, 5388, 5829, -6100, -5085, 6720, 4262, -7243, -3374, 7657, 2432, -7957, -1451, 8135, 445, -8191, 570, 8119, -1580, -7924, 2566, 7603, -3516, -7164, 4412, 6610, -5243, -5952, 5991, 5196, -6647, -4358, 7197, 3446, -7635, -2477, 7949, 1465, -8136, -428, 8190, -620, -8112, 1659, 7897, -2675, -7554, 3647, 7083, -4563, -6494, 5402, 5792, -6155, -4994, 6804, 4107, -7340, -3149, 7751, 2134, -8031, -1081, 8172, 6, -8174, 1071, 8032, -2133, -7750, 3159, 7331, -4133, -6782, 5034, 6110, -5851, -5330, 6562, 4451, -7160, -3491, 7627, 2464, -7960, -1392, 8147, 290, -8187, 818, 8075, -1915, -7816, 2978, 7409, -3989, -6866, 4927, 6190, -5776, -5399, 6516, 4502, -7137, -3520, 7621, 2466, -7963, -1364, 8151, 232, -8185, 905, 8058, -2029, -7775, 3114, 7339, -4142, -6759, 5090, 6043, -5941, -5208, 6674, 4265, -7277, -3237, 7734, 2139, -8039, -999, 8180, -167, -8157, 1330, 7966, -2470, -7613, 3560, 7102, -4581, -6444, 5508, 5649, -6324, -4737, 7007, 3722, -7548, -2628, 7928, 1474, -8144, -289, 8185, -907, -8053, 2084, 7747, -3221, -7275, 4289, 6643, -5268, -5868, 6133, 4961, -6867, -3945, 7451, 2839, -7873, -1669, 8121, 458, -8190, 763, 8075, -1973, -7780, 3138, 7308, -4237, -6672, 5241, 5881, -6129, -4957, 6877, 3915, -7471, -2783, 7893, 1582, -8134, -344, 8186, -906, -8048, 2135, 7720, -3320, -7212, 4426, 6531, -5432, -5695, 6309, 4720, -7039, -3633, 7600, 2454, -7982, -1216, 8170, -57, -8162, 1328, 7954, -2572, -7553, 3753, 6963, -4846, -6204, 5820, 5287, -6654, -4239, 7321, 3082, -7810, -1847, 8101, 561, -8191, 740, 8072, -2026, -7750, 3261, 7229, -4418, -6523, 5461, 5646, -6368, -4624, 7111, 3479, -7672, -2243, 8033, 944, -8187, 381, 8124, -1700, -7849, 2974, 7364, -4174, -6685, 5264, 5824, -6217, -4808, 7003, 3659, -7604, -2411, 8000, 1093)        
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L21C31_i
    );

    L21C32_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-8189, -444, 8116, 1755, -7833, -3020, 7345, 4202, -6670, -5276, 5822, 6209, -4828, -6983, 3710, 7575, -2502, -7975, 1230, 8170, 68, -8160, -1364, 7943, 2621, -7529, -3812, 6926, 4904, -6154, -5874, 5230, 6695, -4180, -7351, 3027, 7824, -1805, -8107, 539, 8190, 735, -8076, -1991, 7766, 3195, -7272, -4321, 6603, 5340, -5780, -6232, 4820, 6973, -3749, -7549, 2591, 7945, -1376, -8157, 129, 8176, 1116, -8007, -2335, 7651, 3495, -7122, -4575, 6429, 5546, -5593, -6390, 4629, 7086, -3564, -7622, 2420, 7984, -1225, -8168, 4, 8168, 1213, -7988, -2403, 7630, 3535, -7107, -4588, 6427, 5538, -5610, -6366, 4671, 7053, -3635, -7588, 2521, 7957, -1356, -8156, 164, 8179, 1028, -8030, -2197, 7710, 3315, -7230, -4364, 6598, 5316, -5832, -6158, 4943, 6869, -3957, -7438, 2889, 7851, -1767, -8105, 608, 8190, 558, -8112, -1712, 7868, 2827, -7468, -3885, 6918, 4862, -6233, -5741, 5424, 6503, -4512, -7137, 3511, 7627, -2446, -7970, 1333, 8154, -199, -8183, -938, 8052, 2053, -7769, -3128, 7336, 4139, -6767, -5071, 6069, 5903, -5260, -6625, 4353, 7219, -3369, -7679, 2322, 7994, -1237, -8163, 129, 8179, 976, -8049, -2063, 7770, 3108, -7353, -4096, 6802, 5007, -6133, -5828, 5354, 6541, -4484, -7138, 3535, 7607, -2527, -7942, 1476, 8136, -403, -8190, -676, 8101, 1738, -7874, -2771, 7510, 3751, -7022, -4668, 6413, 5501, -5699, -6241, 4890, 6873, -4002, -7391, 3049, 7782, -2048, -8046, 1015, 8176, 30, -8173, -1075, 8035, 2097, -7769, -3085, 7376, 4019, -6869, -4889, 6251, 5676, -5537, -6373, 4735, 6967, -3863, -7451, 2930, 7816, -1957, -8061, 953, 8178, 60, -8172, -1072, 8038, 2064, -7785, -3023, 7412, 3932, -6931, -4782, 6345, 5557, -5668, -6248, 4907, 6844, -4077, -7339, 3188, 7723, -2256, -7996, 1292, 8151, -314, -8190, -668, 8109, 1636, -7914, -2580, 7606, 3484, -7194, -4337, 6679, 5126, -6075, -5843, 5386, 6476, -4627, -7020, 3803, 7464, -2933, -7807, 2022, 8041, -1089, -8168, 142, 8184, 803, -8092, -1737, 7891, 2642, -7589, -3513, 7186, 4334, -6692, -5097, 6111, 5791, -5455, -6410, 4729, 6944, -3946, -7390, 3113, 7739, -2246, -7991, 1350, 8141, -442, -8191, -470, 8138, 1372, -7987, -2257, 7737, 3110, -7395, -3925, 6963, 4688, -6450, -5394, 5860, 6033, -5204, -6600, 4486, 7085, -3720, -7489, 2910, 7802, -2071, -8025, 1209, 8154, -337, -8191, -538, 8133, 1403, -7985, -2251, 7745, 3069, -7422, -3853, 7015, 4590, -6534, -5276, 5981, 5900, -5367, -6460, 4693, 6947, -3974, -7359, 3212, 7690, -2420, -7940, 1603, 8104, -774, -8184, -63, 8176, 895, -8086, -1717, 7911, 2517, -7658, -3290, 7326, 4026, -6922, -4721, 6449, 5365, -5915, -5955, 5321, 6483, -4679, -6947, 3992, 7340, -3270, -7662, 2516, 7908, -1743, -8080, 954, 8172, -160, -8188, -635, 8126, 1419, -7990, -2190, 7778, 2936, -7498, -3654, 7148, 4335, -6736, -4976, 6263, 5568, -5737, -6111, 5160, 6596, -4541, -7023, 3883, 7385, -3195, -7684, 2479, 7913, -1747, -8075, 1000, 8167, -249, -8191, -504, 8143, 1247, -8031, -1980, 7850, 2692, -7607, -3381, 7300, 4038, -6938, -4663, 6519, 5245, -6051, -5786, 5535, 6277, -4978, -6719, 4383, 7105, -3758, -7437, 3104, 7708, -2431, -7921, 1739, 8072, -1039, -8163, 332, 8190, 373, -8159, -1075, 8066, 1765, -7916, -2441, 7708, 3095, -7446, -3726, 7130, 4327, -6767, -4896, 6356, 5427, -5903, -5920, 5410, 6369, -4883, -6774, 4322, 7129, -3736, -7437, 3126, 7692, -2499, -7896, 1856, 8046, -1205, -8145, 546, 8188, 111, -8180, -767, 8117, 1413, -8006, -2050, 7842, 2670, -7633, -3272, 7374, 3850, -7074, -4404, 6729, 4927, -6347, -5421, 5927, 5877, -5475, -6299, 4990, 6681, -4480, -7024, 3945, 7322, -3391, -7580, 2817, 7791, -2232, -7960, 1636, 8081, -1034, -8159, 427, 8190, 177, -8177, -780, 8119, 1374, -8020, -1960, 7876, 2532, -7694, -3089, 7470, 3626, -7210, -4144, 6912, 4637, -6583, -5106, 6220, 5545, -5830, -5957, 5410, 6335, -4968, -6683, 4501, 6995, -4017, -7274, 3514, 7515, -2998, -7721, 2469, 7889, -1933, -8021, 1389, 8114, -842, -8172, 293, 8190, 254, -8175, -798, 8121, 1335, -8033, -1865, 7910, 2383, -7755, -2890, 7566, 3380, -7348, -3856, 7099, 4311, -6823, -4749, 6519, 5163, -6192, -5556, 5840, 5923, -5469, -6267, 5076, 6583, -4667, -6874, 4240, 7135, -3801, -7369, 3349, 7573, -2888, -7750, 2417, 7895, -1941, -8013, 1459, 8099, -976, -8159, 491, 8187, -8, -8188, -474, 8159, 950, -8105, -1423, 8022, 1886, -7914, -2342, 7779, 2786, -7621, -3220, 7437, 3640, -7233, -4048, 7005, 4438, -6758, -4815, 6490, 5173, -6206, -5516, 5902, 5837, -5585, -6142, 5251, 6425, -4906, -6689, 4547, 6931, -4179, -7154, 3799, 7354, -3413, -7534, 3018, 7690, -2619, -7827, 2214, 7940, -1807, -8033, 1396, 8103, -986, -8154, 574, 8182, -165, -8191, -244, 8178, 648, -8147, -1049, 8095, 1443, -8026, -1834, 7936, 2215, -7831, -2591, 7706, 2957, -7567, -3315, 7410, 3662, -7239, -4001, 7053, 4326, -6854, -4643, 6640, 4945, -6416, -5237, 6178, 5514, -5932, -5781, 5673, 6032, -5407, -6271, 5131, 6495, -4848, -6707, 4557, 6902, -4261, -7086, 3958, 7253, -3651, -7408, 3339, 7547, -3025, -7674, 2706, 7784, -2387, -7883, 2065, 7966, -1743, -8037, 1420, 8093, -1098, -8138, 776, 8167, -456, -8186, 137, 8190, 178, -8185, -492, 8165, 801, -8136, -1108, 8093, 1409, -8042, -1708, 7978, 1999, -7906, -2288, 7822, 2569, -7731, -2846, 7629, 3115, -7520, -3380, 7401, 3637, -7276, -3888, 7141, 4131, -7002, -4369, 6854, 4598, -6701, -4822, 6541, 5036, -6377, -5245, 6206, 5444, -6032, -5638, 5852, 5822, -5670, -6000, 5482, 6169, -5293, -6333, 5098, 6486, -4903, -6635, 4704, 6774, -4505, -6907, 4302, 7031, -4099, -7150, 3893, 7260, -3689, -7365, 3482, 7461, -3276, -7552, 3068, 7635, -2863, -7713, 2655, 7782, -2451, -7848, 2245, 7905, -2042, -7958, 1838, 8004, -1638, -8046, 1437, 8080, -1240, -8112, 1043, 8136, -849, -8157, 656, 8171, -467, -8183, 278, 8188, -94, -8191, -90, 8189, 269, -8184, -448, 8173, 622, -8161, -794, 8143, 962, -8124, -1129, 8101, 1291, -8076, -1452, 8046, 1608, -8016, -1762, 7982, 1912, -7947, -2060, 7908, 2203, -7869, -2345, 7827, 2481, -7785, -2617, 7739, 2747, -7694, -2876, 7645, 3000, -7598, -3122, 7547, 3240, -7498, -3356, 7446, 3467, -7395, -3577, 7342, 3682, -7291, -3786, 7237, 3885, -7185, -3983, 7131, 4076, -7079, -4167, 7025, 4255, -6973, -4341, 6920, 4422, -6869, -4503, 6817, 4578, -6767, -4654, 6716, 4724, -6667, -4794, 6617, 4859, -6570, -4924, 6523, 4984, -6478, -5043, 6432, 5099, -6389, -5154, 6345, 5204, -6305, -5254, 6264, 5300, -6226, -5346, 6188, 5387, -6153, -5428, 6117, 5465, -6085, -5502, 6052, 5535, -6023, -5568, 5994, 5596, -5968, -5625, 5942, 5650, -5919, -5674, 5896, 5695, -5877, -5716, 5858, 5733, -5842, -5750, 5826, 5763, -5814, -5776, 5802, 5786, -5794, -5795, 5785, 5801, -5780, -5807, 5775, 5809, -5774, -5811, 5772, 5810, -5775, -5808, 5777, 5803, -5783, -5798, 5789, 5789, -5799, -5781, 5809, 5768, -5822, -5756, 5835, 5739, -5852, -5723, 5869, 5703, -5890, -5683, 5910, 5659, -5934, -5635, 5957, 5607, -5984, -5579, 6011, 5547, -6042, -5515, 6072, 5479, -6105, -5443, 6138, 5402, -6175, -5362, 6211, 5317, -6250, -5272, 6289, 5223, -6331, -5173, 6372, 5119, -6416, -5065, 6459, 5006, -6506, -4947, 6552, 4883, -6600, -4819, 6647, 4750, -6698, -4681, 6747, 4607, -6798, -4532, 6849, 4453, -6901, -4372, 6952, 4287, -7006, -4201, 7058, 4110, -7112, -4019, 7164, 3922, -7218, -3824, 7270, 3721, -7323, -3618, 7375, 3509, -7428, -3399, 7478, 3284, -7529, -3168, 7578, 3046, -7628, -2924, 7675, 2796, -7723, -2667, 7767, 2533, -7812, -2397, 7853, 2257, -7894, -2115, 7932, 1968, -7969, -1820, 8003, 1666, -8036, -1512, 8064, 1352, -8092, -1191, 8115, 1026, -8137, -859, 8154, 687, -8169, -514, 8179, 337, -8188, -159, 8190, -24, -8191, 207, 8185, -395, -8177, 583, 8162, -776, -8145, 969, 8121, -1165, -8093, 1362, 8059, -1562, -8021, 1762, 7976, -1965, -7927, 2168, 7870, -2373, -7809, 2578, 7739, -2785, -7666, 2990, 7584, -3198, -7497, 3403, 7402, -3611, -7302, 3816, 7192, -4022, -7078, 4225, 6955, -4428, -6826, 4628, 6688, -4829, -6544, 5024, 6391, -5220, -6233, 5410, 6065, -5599, -5891, 5783, 5708, -5965, -5519, 6140, 5320, -6313, -5116, 6479, 4903, -6642, -4684, 6796, 4456, -6947, -4223, 7089, 3981, -7226, -3733, 7354, 3478, -7476, -3217, 7588, 2948, -7694, -2675, 7788, 2394, -7876, -2110, 7951, 1818, -8019, -1523, 8075, 1222, -8121, -918, 8155, 609, -8179, -298, 8189, -18, -8190, 334, 8176, -655, -8151, 975, 8111, -1298, -8060, 1620, 7994, -1944, -7917, 2265, 7823, -2586, -7718, 2904, 7596, -3221, -7463, 3533, 7313, -3843, -7151, 4146, 6973, -4446, -6783, 4738, 6576, -5025, -6358, 5303, 6124, -5574, -5878, 5834, 5616, -6087, -5344, 6327, 5057, -6557, -4759, 6774, 4447, -6979, -4126, 7170, 3791, -7348, -3448, 7509, 3093, -7656, -2731, 7785, 2358, -7899, -1979, 7993, 1592, -8072, -1199, 8129, 800, -8170, -398, 8188, -10, -8189, 418, 8167, -830, -8126, 1240, 8062, -1652, -7978, 2060, 7872, -2466, -7745, 2867, 7595, -3265, -7425, 3653, 7232, -4036, -7019, 4408, 6783, -4772, -6528, 5122, 6251, -5461, -5956, 5784, 5639, -6093, -5306, 6384, 4952, -6659, -4584, 6913, 4197, -7149, -3797, 7362, 3380, -7554, -2952, 7721, 2510, -7866, -2060, 7983, 1598, -8077, -1131, 8142, 655, -8181, -176, 8190, -308, -8173, 792, 8125, -1277, -8050, 1758, 7943, -2238, -7809, 2710, 7643, -3176, -7450, 3631, 7227, -4076, -6976, 4506, 6696, -4923, -6390, 5321, 6056, -5702, -5699, 6061, 5314, -6399, -4909, 6710, 4479, -6998, -4031, 7256, 3562, -7488, -3078, 7687, 2576, -7856, -2063, 7990, 1536, -8092, -1003, 8158, 460, -8189, 85, 8183, -634, -8141, 1182, 8060, -1728, -7944, 2267, 7789, -2800, -7598, 3320, 7369, -3829, -7105, 4319, 6804, -4794, -6471, 5245, 6103, -5674, -5705, 6075, 5275, -6450, -4818, 6791, 4333, -7102, -3826, 7375, 3294, -7614, -2745, 7811, 2178, -7971, -1598, 8086, 1005, -8161, -407, 8190, -199, -8176, 804, 8115, -1409, -8011, 2007, 7860, -2598, -7666, 3175, 7425, -3738, -7142, 4279, 6815, -4801, -6449, 5294, 6041, -5760, -5598, 6191, 5118, -6589, -4606, 6947, 4063, -7266, -3495, 7539, 2900, -7769, -2287, 7949, 1656, -8082, -1013, 8162, 360, -8191, 297, 8166, -956, -8090, 1610, 7959, -2257, -7776, 2890, 7539, -3508, -7252, 4103, 6914, -4674, -6528, 5213, 6095, -5721, -5619, 6189, 5101, -6617, -4547, 6998, 3957, -7333, -3338, 7615, 2691, -7844, -2024, 8016, 1337, -8131, -641, 8185, -65, -8181, 771, 8113, -1476, -7986, 2170, 7795, -2852, -7547, 3513, 7237, -4151, -6872, 4756, 6451, -5329, -5978, 5860, 5455, -6348, -4889, 6785, 4279, -7170, -3634, 7497, 2956, -7766, -2252, 7969, 1526, -8109, -787, 8180, 36, -8184, 715, 8118, -1465, -7983, 2203, 7778, -2927, -7506, 3625, 7167, -4296, -6765, 4930, 6301, -5525, -5781, 6070, 5206, -6564, -4584, 6999, 3916, -7373, -3212, 7680, 2475, -7918, -1714, 8083, 933, -8174, -142, 8187, -654, -8124, 1445, 7982, -2226, -7765, 2987, 7470, -3723, -7104, 4423, 6666, -5084, -6163, 5696, 5595, -6254, -4972, 6750, 4294, -7182, -3574, 7540, 2813, -7825, -2023, 8029, 1208, -8153, -380, 8190, -457, -8145, 1290, 8011, -2113, -7795, 2915, 7493, -3690, -7113, 4426, 6652, -5118, -6121, 5755, 5519, -6333, -4857, 6841, 4137, -7278, -3371, 7632, 2564, -7905, -1727, 8087, 867, -8180, 4, 8179, -880, -8085, 1746, 7897, -2596, -7618, 3417, 7248, -4202, -6794, 4938, 6256, -5620, -5645, 6235, 4962, -6779, -4221, 7241, 3424, -7619, -2585, 7903, 1710, -8093, -814, 8183, -97, -8173, 1007, 8059, -1909, -7847, 2788, 7532, -3636, -7124, 4438, 6622, -5188, -6036, 5871, 5368, -6482, -4631, 7009, 3830, -7448, -2978, 7788, 2083, -8029, -1160, 8161, 216, -8187, 730, 8102, -1672, -7908, 2591, 7605, -3479, -7200, 4321, 6693, -5107, -6094, 5823, 5407, -6462, -4645, 7010, 3813, -7463, -2928, 7810, 1997, -8049, -1037, 8172, 58, -8180, 922, 8068, -1894, -7841, 2839, 7497, -3747, -7044, 4600, 6485, -5389, -5830, 6099, 5084, -6721, -4263, 7242, 3373, -7658, -2433, 7956, 1450, -8136, -446, 8190, -571, -8120, 1579, 7923, -2567, -7604, 3515, 7163, -4413, -6611, 5242, 5951, -5992, -5197, 6646, 4357, -7198, -3447, 7634, 2476, -7950, -1466, 8135, 427, -8191, 619, 8111, -1660, -7898, 2674, 7553, -3648, -7084, 4562, 6493, -5403, -5793, 6154, 4993, -6805, -4108, 7339, 3148, -7752, -2135, 8030, 1080, -8173, -7, 8173, -1072, -8033, 2132, 7749, -3160, -7332, 4132, 6781, -5035, -6111, 5850, 5329, -6563, -4452, 7159, 3490, -7628, -2465, 7959, 1391, -8148, -291, 8186, -819, -8076, 1914, 7815, -2979, -7410, 3988, 6865, -4928, -6191, 5775, 5398, -6517, -4503, 7136, 3519, -7622, -2467, 7962, 1363, -8152, -233, 8184, -906, -8059, 2028, 7774, -3115, -7340, 4141, 6758, -5091, -6044, 5940, 5207, -6675, -4266, 7276, 3236, -7735, -2140, 8038, 998, -8181, 166, 8156, -1331, -7967, 2469, 7612, -3561, -7103, 4580, 6443, -5509, -5650, 6323, 4736, -7008, -3723, 7547, 2627, -7929, -1475, 8143, 288, -8186, 906, 8052, -2085, -7748, 3220, 7274, -4290, -6644, 5267, 5867, -6134, -4962, 6866, 3944, -7452, -2840, 7872, 1668, -8122, -459, 8189, -764, -8076, 1972, 7779, -3139, -7309, 4236, 6671, -5242, -5882, 6128, 4956, -6878, -3916, 7470, 2782, -7894, -1583, 8133, 343, -8187, 905, 8047, -2136, -7721, 3319, 7211, -4427, -6532, 5431, 5694, -6310, -4721, 7038, 3632, -7601, -2455, 7981, 1215, -8171, 56, 8161, -1329, -7955, 2571, 7552, -3754, -6964, 4845, 6203, -5821, -5288, 6653, 4238, -7322, -3083, 7809, 1846, -8102, -562, 8190, -741, -8073, 2025, 7749, -3262, -7230, 4417, 6522, -5462, -5647, 6367, 4623, -7112, -3480, 7671, 2242, -8034, -945, 8186, -382, -8125, 1699, 7848, -2975, -7365, 4173, 6684, -5265, -5825, 6216, 4807, -7004, -3660, 7603, 2410, -8001, -1094)    
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L21C32_i
    );

    L21C33_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (8188, 443, -8117, -1756, 7832, 3019, -7346, -4203, 6669, 5275, -5823, -6210, 4827, 6982, -3711, -7576, 2501, 7974, -1231, -8171, -69, 8159, 1363, -7944, -2622, 7528, 3811, -6927, -4905, 6153, 5873, -5231, -6696, 4179, 7350, -3028, -7825, 1804, 8106, -540, -8191, -736, 8075, 1990, -7767, -3196, 7271, 4320, -6604, -5341, 5779, 6231, -4821, -6974, 3748, 7548, -2592, -7946, 1375, 8156, -130, -8177, -1117, 8006, 2334, -7652, -3496, 7121, 4574, -6430, -5547, 5592, 6389, -4630, -7087, 3563, 7621, -2421, -7985, 1224, 8167, -5, -8169, -1214, 7987, 2402, -7631, -3536, 7106, 4587, -6428, -5539, 5609, 6365, -4672, -7054, 3634, 7587, -2522, -7958, 1355, 8155, -165, -8180, -1029, 8029, 2196, -7711, -3316, 7229, 4363, -6599, -5317, 5831, 6157, -4944, -6870, 3956, 7437, -2890, -7852, 1766, 8104, -609, -8191, -559, 8111, 1711, -7869, -2828, 7467, 3884, -6919, -4863, 6232, 5740, -5425, -6504, 4511, 7136, -3512, -7628, 2445, 7969, -1334, -8155, 198, 8182, 937, -8053, -2054, 7768, 3127, -7337, -4140, 6766, 5070, -6070, -5904, 5259, 6624, -4354, -7220, 3368, 7678, -2323, -7995, 1236, 8162, -130, -8180, -977, 8048, 2062, -7771, -3109, 7352, 4095, -6803, -5008, 6132, 5827, -5355, -6542, 4483, 7137, -3536, -7608, 2526, 7941, -1477, -8137, 402, 8189, 675, -8102, -1739, 7873, 2770, -7511, -3752, 7021, 4667, -6414, -5502, 5698, 6240, -4891, -6874, 4001, 7390, -3050, -7783, 2047, 8045, -1016, -8177, -31, 8172, 1074, -8036, -2098, 7768, 3084, -7377, -4020, 6868, 4888, -6252, -5677, 5536, 6372, -4736, -6968, 3862, 7450, -2931, -7817, 1956, 8060, -954, -8179, -61, 8171, 1071, -8039, -2065, 7784, 3022, -7413, -3933, 6930, 4781, -6346, -5558, 5667, 6247, -4908, -6845, 4076, 7338, -3189, -7724, 2255, 7995, -1293, -8152, 313, 8189, 667, -8110, -1637, 7913, 2579, -7607, -3485, 7193, 4336, -6680, -5127, 6074, 5842, -5387, -6477, 4626, 7019, -3804, -7465, 2932, 7806, -2023, -8042, 1088, 8167, -143, -8185, -804, 8091, 1736, -7892, -2643, 7588, 3512, -7187, -4335, 6691, 5096, -6112, -5792, 5454, 6409, -4730, -6945, 3945, 7389, -3114, -7740, 2245, 7990, -1351, -8142, 441, 8190, 469, -8139, -1373, 7986, 2256, -7738, -3111, 7394, 3924, -6964, -4689, 6449, 5393, -5861, -6034, 5203, 6599, -4487, -7086, 3719, 7488, -2911, -7803, 2070, 8024, -1210, -8155, 336, 8190, 537, -8134, -1404, 7984, 2250, -7746, -3070, 7421, 3852, -7016, -4591, 6533, 5275, -5982, -5901, 5366, 6459, -4694, -6948, 3973, 7358, -3213, -7691, 2419, 7939, -1604, -8105, 773, 8183, 62, -8177, -896, 8085, 1716, -7912, -2518, 7657, 3289, -7327, -4027, 6921, 4720, -6450, -5366, 5914, 5954, -5322, -6484, 4678, 6946, -3993, -7341, 3269, 7661, -2517, -7909, 1742, 8079, -955, -8173, 159, 8187, 634, -8127, -1420, 7989, 2189, -7779, -2937, 7497, 3653, -7149, -4336, 6735, 4975, -6264, -5569, 5736, 6110, -5161, -6597, 4540, 7022, -3884, -7386, 3194, 7683, -2480, -7914, 1746, 8074, -1001, -8168, 248, 8190, 503, -8144, -1248, 8030, 1979, -7851, -2693, 7606, 3380, -7301, -4039, 6937, 4662, -6520, -5246, 6050, 5785, -5536, -6278, 4977, 6718, -4384, -7106, 3757, 7436, -3105, -7709, 2430, 7920, -1740, -8073, 1038, 8162, -333, -8191, -374, 8158, 1074, -8067, -1766, 7915, 2440, -7709, -3096, 7445, 3725, -7131, -4328, 6766, 4895, -6357, -5428, 5902, 5919, -5411, -6370, 4882, 6773, -4323, -7130, 3735, 7436, -3127, -7693, 2498, 7895, -1857, -8047, 1204, 8144, -547, -8189, -112, 8179, 766, -8118, -1414, 8005, 2049, -7843, -2671, 7632, 3271, -7375, -3851, 7073, 4403, -6730, -4928, 6346, 5420, -5928, -5878, 5474, 6298, -4991, -6682, 4479, 7023, -3946, -7323, 3390, 7579, -2818, -7792, 2231, 7959, -1637, -8082, 1033, 8158, -428, -8191, -178, 8176, 779, -8120, -1375, 8019, 1959, -7877, -2533, 7693, 3088, -7471, -3627, 7209, 4143, -6913, -4638, 6582, 5105, -6221, -5546, 5829, 5956, -5411, -6336, 4967, 6682, -4502, -6996, 4016, 7273, -3515, -7516, 2997, 7720, -2470, -7890, 1932, 8020, -1390, -8115, 841, 8171, -294, -8191, -255, 8174, 797, -8122, -1336, 8032, 1864, -7911, -2384, 7754, 2889, -7567, -3381, 7347, 3855, -7100, -4312, 6822, 4748, -6520, -5164, 6191, 5555, -5841, -5924, 5468, 6266, -5077, -6584, 4666, 6873, -4241, -7136, 3800, 7368, -3350, -7574, 2887, 7749, -2418, -7896, 1940, 8012, -1460, -8100, 975, 8158, -492, -8188, 7, 8187, 473, -8160, -951, 8104, 1422, -8023, -1887, 7913, 2341, -7780, -2787, 7620, 3219, -7438, -3641, 7232, 4047, -7006, -4439, 6757, 4814, -6491, -5174, 6205, 5515, -5903, -5838, 5584, 6141, -5252, -6426, 4905, 6688, -4548, -6932, 4178, 7153, -3800, -7355, 3412, 7533, -3019, -7691, 2618, 7826, -2215, -7941, 1806, 8032, -1397, -8104, 985, 8153, -575, -8183, 164, 8190, 243, -8179, -649, 8146, 1048, -8096, -1444, 8025, 1833, -7937, -2216, 7830, 2590, -7707, -2958, 7566, 3314, -7411, -3663, 7238, 4000, -7054, -4327, 6853, 4642, -6641, -4946, 6415, 5236, -6179, -5515, 5931, 5780, -5674, -6033, 5406, 6270, -5132, -6496, 4847, 6706, -4558, -6903, 4260, 7085, -3959, -7254, 3650, 7407, -3340, -7548, 3024, 7673, -2707, -7785, 2386, 7882, -2066, -7967, 1742, 8036, -1421, -8094, 1097, 8137, -777, -8168, 455, 8185, -138, -8191, -179, 8184, 491, -8166, -802, 8135, 1107, -8094, -1410, 8041, 1707, -7979, -2000, 7905, 2287, -7823, -2570, 7730, 2845, -7630, -3116, 7519, 3379, -7402, -3638, 7275, 3887, -7142, -4132, 7001, 4368, -6855, -4599, 6700, 4821, -6542, -5037, 6376, 5244, -6207, -5445, 6031, 5637, -5853, -5823, 5669, 5999, -5483, -6170, 5292, 6332, -5099, -6487, 4902, 6634, -4705, -6775, 4504, 6906, -4303, -7032, 4098, 7149, -3894, -7261, 3688, 7364, -3483, -7462, 3275, 7551, -3069, -7636, 2862, 7712, -2656, -7783, 2450, 7847, -2246, -7906, 2041, 7957, -1839, -8005, 1637, 8045, -1438, -8081, 1239, 8111, -1044, -8137, 848, 8156, -657, -8172, 466, 8182, -279, -8189, 93, 8190, 89, -8190, -270, 8183, 447, -8174, -623, 8160, 793, -8144, -963, 8123, 1128, -8102, -1292, 8075, 1451, -8047, -1609, 8015, 1761, -7983, -1913, 7946, 2059, -7909, -2204, 7868, 2344, -7828, -2482, 7784, 2616, -7740, -2748, 7693, 2875, -7646, -3001, 7597, 3121, -7548, -3241, 7497, 3355, -7447, -3468, 7394, 3576, -7343, -3683, 7290, 3785, -7238, -3886, 7184, 3982, -7132, -4077, 7078, 4166, -7026, -4256, 6972, 4340, -6921, -4423, 6868, 4502, -6818, -4579, 6766, 4653, -6717, -4725, 6666, 4793, -6618, -4860, 6569, 4923, -6524, -4985, 6477, 5042, -6433, -5100, 6388, 5153, -6346, -5205, 6304, 5253, -6265, -5301, 6225, 5345, -6189, -5388, 6152, 5427, -6118, -5466, 6084, 5501, -6053, -5536, 6022, 5567, -5995, -5597, 5967, 5624, -5943, -5651, 5918, 5673, -5897, -5696, 5876, 5715, -5859, -5734, 5841, 5749, -5827, -5764, 5813, 5775, -5803, -5787, 5793, 5794, -5786, -5802, 5779, 5806, -5776, -5810, 5773, 5810, -5773, -5811, 5774, 5807, -5778, -5804, 5782, 5797, -5790, -5790, 5798, 5780, -5810, -5769, 5821, 5755, -5836, -5740, 5851, 5722, -5870, -5704, 5889, 5682, -5911, -5660, 5933, 5634, -5958, -5608, 5983, 5578, -6012, -5548, 6041, 5514, -6073, -5480, 6104, 5442, -6139, -5403, 6174, 5361, -6212, -5318, 6249, 5271, -6290, -5224, 6330, 5172, -6373, -5120, 6415, 5064, -6460, -5007, 6505, 4946, -6553, -4884, 6599, 4818, -6648, -4751, 6697, 4680, -6748, -4608, 6797, 4531, -6850, -4454, 6900, 4371, -6953, -4288, 7005, 4200, -7059, -4111, 7111, 4018, -7165, -3923, 7217, 3823, -7271, -3722, 7322, 3617, -7376, -3510, 7427, 3398, -7479, -3285, 7528, 3167, -7579, -3047, 7627, 2923, -7676, -2797, 7722, 2666, -7768, -2534, 7811, 2396, -7854, -2258, 7893, 2114, -7933, -1969, 7968, 1819, -8004, -1667, 8035, 1511, -8065, -1353, 8091, 1190, -8116, -1027, 8136, 858, -8155, -688, 8168, 513, -8180, -338, 8187, 158, -8191, 23, 8190, -208, -8186, 394, 8176, -584, -8163, 775, 8144, -970, -8122, 1164, 8092, -1363, -8060, 1561, 8020, -1763, -7977, 1964, 7926, -2169, -7871, 2372, 7808, -2579, -7740, 2784, 7665, -2991, -7585, 3197, 7496, -3404, -7403, 3610, 7301, -3817, -7193, 4021, 7077, -4226, -6956, 4427, 6825, -4629, -6689, 4828, 6543, -5025, -6392, 5219, 6232, -5411, -6066, 5598, 5890, -5784, -5709, 5964, 5518, -6141, -5321, 6312, 5115, -6480, -4904, 6641, 4683, -6797, -4457, 6946, 4222, -7090, -3982, 7225, 3732, -7355, -3479, 7475, 3216, -7589, -2949, 7693, 2674, -7789, -2395, 7875, 2109, -7952, -1819, 8018, 1522, -8076, -1223, 8120, 917, -8156, -610, 8178, 297, -8190, 17, 8189, -335, -8177, 654, 8150, -976, -8112, 1297, 8059, -1621, -7995, 1943, 7916, -2266, -7824, 2585, 7717, -2905, -7597, 3220, 7462, -3534, -7314, 3842, 7150, -4147, -6974, 4445, 6782, -4739, -6577, 5024, 6357, -5304, -6125, 5573, 5877, -5835, -5617, 6086, 5343, -6328, -5058, 6556, 4758, -6775, -4448, 6978, 4125, -7171, -3792, 7347, 3447, -7510, -3094, 7655, 2730, -7786, -2359, 7898, 1978, -7994, -1593, 8071, 1198, -8130, -801, 8169, 397, -8189, 9, 8188, -419, -8168, 829, 8125, -1241, -8063, 1651, 7977, -2061, -7873, 2465, 7744, -2868, -7596, 3264, 7424, -3654, -7233, 4035, 7018, -4409, -6784, 4771, 6527, -5123, -6252, 5460, 5955, -5785, -5640, 6092, 5305, -6385, -4953, 6658, 4583, -6914, -4198, 7148, 3796, -7363, -3381, 7553, 2951, -7722, -2511, 7865, 2059, -7984, -1599, 8076, 1130, -8143, -656, 8180, 175, -8191, 307, 8172, -793, -8126, 1276, 8049, -1759, -7944, 2237, 7808, -2711, -7644, 3175, 7449, -3632, -7228, 4075, 6975, -4507, -6697, 4922, 6389, -5322, -6057, 5701, 5698, -6062, -5315, 6398, 4908, -6711, -4480, 6997, 4030, -7257, -3563, 7487, 3077, -7688, -2577, 7855, 2062, -7991, -1537, 8091, 1002, -8159, -461, 8188, -86, -8184, 633, 8140, -1183, -8061, 1727, 7943, -2268, -7790, 2799, 7597, -3321, -7370, 3828, 7104, -4320, -6805, 4793, 6470, -5246, -6104, 5673, 5704, -6076, -5276, 6449, 4817, -6792, -4334, 7101, 3825, -7376, -3295, 7613, 2744, -7812, -2179, 7970, 1597, -8087, -1006, 8160, 406, -8191, 198, 8175, -805, -8116, 1408, 8010, -2008, -7861, 2597, 7665, -3176, -7426, 3737, 7141, -4280, -6816, 4800, 6448, -5295, -6042, 5759, 5597, -6192, -5119, 6588, 4605, -6948, -4064, 7265, 3494, -7540, -2901, 7768, 2286, -7950, -1657, 8081, 1012, -8163, -361, 8190, -298, -8167, 955, 8089, -1611, -7960, 2256, 7775, -2891, -7540, 3507, 7251, -4104, -6915, 4673, 6527, -5214, -6096, 5720, 5618, -6190, -5102, 6616, 4546, -6999, -3958, 7332, 3337, -7616, -2692, 7843, 2023, -8017, -1338, 8130, 640, -8186, 64, 8180, -772, -8114, 1475, 7985, -2171, -7796, 2851, 7546, -3514, -7238, 4150, 6871, -4757, -6452, 5328, 5977, -5861, -5456, 6347, 4888, -6786, -4280, 7169, 3633, -7498, -2957, 7765, 2251, -7970, -1527, 8108, 786, -8181, -37, 8183, -716, -8119, 1464, 7982, -2204, -7779, 2926, 7505, -3626, -7168, 4295, 6764, -4931, -6302, 5524, 5780, -6071, -5207, 6563, 4583, -7000, -3917, 7372, 3211, -7681, -2476, 7917, 1713, -8084, -934, 8173, 141, -8188, 653, 8123, -1446, -7983, 2225, 7764, -2988, -7471, 3722, 7103, -4424, -6667, 5083, 6162, -5697, -5596, 6253, 4971, -6751, -4295, 7181, 3573, -7541, -2814, 7824, 2022, -8030, -1209, 8152, 379, -8191, 456, 8144, -1291, -8012, 2112, 7794, -2916, -7494, 3689, 7112, -4427, -6653, 5117, 6120, -5756, -5520, 6332, 4856, -6842, -4138, 7277, 3370, -7633, -2565, 7904, 1726, -8088, -868, 8179, -5, -8180, 879, 8084, -1747, -7898, 2595, 7617, -3418, -7249, 4201, 6793, -4939, -6257, 5619, 5644, -6236, -4963, 6778, 4220, -7242, -3425, 7618, 2584, -7904, -1711, 8092, 813, -8184, 96, 8172, -1008, -8060, 1908, 7846, -2789, -7533, 3635, 7123, -4439, -6623, 5187, 6035, -5872, -5369, 6481, 4630, -7010, -3831, 7447, 2977, -7789, -2084, 8028, 1159, -8162, -217, 8186, -731, -8103, 1671, 7907, -2592, -7606, 3478, 7199, -4322, -6694, 5106, 6093, -5824, -5408, 6461, 4644, -7011, -3814, 7462, 2927, -7811, -1998, 8048, 1036, -8173, -59, 8179, -923, -8069, 1893, 7840, -2840, -7498, 3746, 7043, -4601, -6486, 5388, 5829, -6100, -5085, 6720, 4262, -7243, -3374, 7657, 2432, -7957, -1451, 8135, 445, -8191, 570, 8119, -1580, -7924, 2566, 7603, -3516, -7164, 4412, 6610, -5243, -5952, 5991, 5196, -6647, -4358, 7197, 3446, -7635, -2477, 7949, 1465, -8136, -428, 8190, -620, -8112, 1659, 7897, -2675, -7554, 3647, 7083, -4563, -6494, 5402, 5792, -6155, -4994, 6804, 4107, -7340, -3149, 7751, 2134, -8031, -1081, 8172, 6, -8174, 1071, 8032, -2133, -7750, 3159, 7331, -4133, -6782, 5034, 6110, -5851, -5330, 6562, 4451, -7160, -3491, 7627, 2464, -7960, -1392, 8147, 290, -8187, 818, 8075, -1915, -7816, 2978, 7409, -3989, -6866, 4927, 6190, -5776, -5399, 6516, 4502, -7137, -3520, 7621, 2466, -7963, -1364, 8151, 232, -8185, 905, 8058, -2029, -7775, 3114, 7339, -4142, -6759, 5090, 6043, -5941, -5208, 6674, 4265, -7277, -3237, 7734, 2139, -8039, -999, 8180, -167, -8157, 1330, 7966, -2470, -7613, 3560, 7102, -4581, -6444, 5508, 5649, -6324, -4737, 7007, 3722, -7548, -2628, 7928, 1474, -8144, -289, 8185, -907, -8053, 2084, 7747, -3221, -7275, 4289, 6643, -5268, -5868, 6133, 4961, -6867, -3945, 7451, 2839, -7873, -1669, 8121, 458, -8190, 763, 8075, -1973, -7780, 3138, 7308, -4237, -6672, 5241, 5881, -6129, -4957, 6877, 3915, -7471, -2783, 7893, 1582, -8134, -344, 8186, -906, -8048, 2135, 7720, -3320, -7212, 4426, 6531, -5432, -5695, 6309, 4720, -7039, -3633, 7600, 2454, -7982, -1216, 8170, -57, -8162, 1328, 7954, -2572, -7553, 3753, 6963, -4846, -6204, 5820, 5287, -6654, -4239, 7321, 3082, -7810, -1847, 8101, 561, -8191, 740, 8072, -2026, -7750, 3261, 7229, -4418, -6523, 5461, 5646, -6368, -4624, 7111, 3479, -7672, -2243, 8033, 944, -8187, 381, 8124, -1700, -7849, 2974, 7364, -4174, -6685, 5264, 5824, -6217, -4808, 7003, 3659, -7604, -2411, 8000, 1093)        
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L21C33_i
    );

    L32_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-2124, -8057, 819, 8189, 504, -8108, -1815, 7815, 3074, -7320, -4254, 6635, 5320, -5780, -6250, 4776, 7015, -3652, -7601, 2434, 7990, -1158, -8176, -149, 8151, 1448, -7921, -2711, 7489, 3901, -6870, -4993, 6076, 5956, -5133, -6770, 4060, 7412, -2889, -7869, 1646, 8128, -365, -8187, -925, 8040, 2189, -7697, -3399, 7163, 4521, -6455, -5533, 5588, 6407, -4587, -7124, 3474, 7665, -2280, -8022, 1030, 8181, 241, -8144, -1506, 7910, 2732, -7487, -3892, 6884, 4956, -6119, -5902, 5208, 6704, -4175, -7348, 3043, 7815, -1843, -8099, 599, 8190, 655, -8091, -1895, 7800, 3086, -7330, -4206, 6687, 5224, -5893, -6122, 4960, 6875, -3917, -7471, 2783, 7892, -1588, -8133, 357, 8186, 879, -8055, -2095, 7738, 3260, -7248, -4351, 6593, 5341, -5792, -6211, 4860, 6938, -3823, -7511, 2699, 7913, -1519, -8140, 304, 8185, 913, -8050, -2110, 7736, 3258, -7253, -4334, 6610, 5311, -5826, -6173, 4913, 6898, -3897, -7473, 2795, 7883, -1637, -8125, 443, 8189, 757, -8079, -1941, 7794, 3080, -7345, -4153, 6738, 5135, -5991, -6008, 5116, 6751, -4136, -7352, 3068, 7796, -1940, -8078, 771, 8189, 411, -8130, -1585, 7901, 2721, -7510, -3802, 6963, 4801, -6275, -5702, 5457, 6482, -4531, -7131, 3511, 7631, -2423, -7978, 1286, 8160, -126, -8179, -1036, 8031, 2174, -7724, -3268, 7260, 4294, -6655, -5234, 5915, 6067, -5062, -6781, 4107, 7357, -3075, -7790, 1982, 8066, -853, -8187, -292, 8145, 1428, -7947, -2537, 7592, 3593, -7094, -4579, 6457, 5474, -5699, -6265, 4831, 6932, -3874, -7468, 2842, 7859, -1760, -8102, 644, 8190, 480, -8125, -1596, 7906, 2677, -7540, -3709, 7032, 4669, -6396, -5542, 5640, 6309, -4783, -6960, 3837, 7479, -2824, -7863, 1759, 8100, -665, -8191, -442, 8130, 1536, -7924, -2603, 7573, 3620, -7089, -4571, 6475, 5438, -5748, -6207, 4918, 6863, -4004, -7397, 3018, 7798, -1982, -8062, 911, 8182, 173, -8160, -1253, 7994, 2309, -7690, -3324, 7251, 4278, -6689, -5158, 6010, 5946, -5231, -6633, 4362, 7203, -3421, -7651, 2421, 7966, -1384, -8147, 323, 8188, 740, -8093, -1790, 7860, 2807, -7498, -3777, 7009, 4681, -6406, -5507, 5696, 6239, -4895, -6869, 4013, 7382, -3068, -7776, 2072, 8040, -1047, -8175, 4, 8174, 1036, -8043, -2059, 7781, 3045, -7396, -3983, 6891, 4853, -6279, -5646, 5566, 6347, -4768, -6948, 3894, 7436, -2962, -7808, 1983, 8055, -976, -8178, -46, 8172, 1063, -8040, -2065, 7783, 3031, -7407, -3950, 6917, 4806, -6324, -5588, 5633, 6282, -4859, -6881, 4011, 7374, -3106, -7756, 2154, 8019, -1174, -8164, 175, 8184, 823, -8085, -1808, 7864, 2764, -7529, -3678, 7082, 4536, -6534, -5327, 5889, 6037, -5162, -6660, 4359, 7184, -3496, -7605, 2583, 7913, -1636, -8110, 665, 8189, 312, -8152, -1284, 7999, 2235, -7734, -3154, 7359, 4025, -6883, -4841, 6310, 5585, -5652, -6252, 4915, 6830, -4112, -7314, 3253, 7694, -2353, -7971, 1419, 8136, -471, -8191, -485, 8134, 1430, -7969, -2356, 7695, 3247, -7320, -4095, 6845, 4884, -6283, -5610, 5636, 6257, -4918, -6823, 4134, 7296, -3299, -7674, 2421, 7950, -1515, -8123, 589, 8190, 341, -8152, -1267, 8007, 2173, -7762, -3052, 7417, 3888, -6979, -4675, 6452, 5399, -5847, -6056, 5167, 6634, -4426, -7130, 3628, 7534, -2790, -7845, 1916, 8057, -1022, -8172, 115, 8184, 789, -8097, -1684, 7911, 2555, -7630, -3395, 7256, 4191, -6797, -4937, 6256, 5620, -5643, -6237, 4962, 6777, -4225, -7237, 3438, 7609, -2614, -7893, 1759, 8083, -887, -8179, 5, 8179, 874, -8086, -1743, 7898, 2589, -7622, -3405, 7257, 4178, -6813, -4905, 6290, 5573, -5699, -6178, 5043, 6711, -4334, -7170, 3576, 7547, -2782, -7840, 1957, 8045, -1113, -8163, 258, 8189, 597, -8127, -1446, 7976, 2275, -7740, -3080, 7419, 3849, -7022, -4576, 6548, 5251, -6007, -5871, 5402, 6426, -4743, -6913, 4033, 7326, -3285, -7662, 2501, 7916, -1696, -8090, 872, 8178, -44, -8183, -786, 8103, 1604, -7942, -2405, 7699, 3179, -7380, -3921, 6986, 4620, -6524, -5273, 5997, 5871, -5413, -6410, 4774, 6884, -4092, -7291, 3369, 7623, -2616, -7882, 1838, 8062, -1046, -8166, 243, 8189, 558, -8135, -1355, 8002, 2135, -7795, -2894, 7513, 3623, -7162, -4318, 6743, 4970, -6264, -5575, 5725, 6125, -5137, -6620, 4501, 7051, -3827, -7418, 3117, 7714, -2382, -7942, 1626, 8096, -858, -8178, 83, 8185, 690, -8121, -1457, 7983, 2207, -7776, -2938, 7500, 3639, -7160, -4309, 6757, 4938, -6298, -5525, 5784, 6061, -5223, -6546, 4616, 6971, -3974, -7339, 3297, 7641, -2596, -7880, 1873, 8051, -1138, -8156, 393, 8190, 352, -8159, -1094, 8059, 1823, -7895, -2538, 7665, 3228, -7375, -3893, 7025, 4522, -6620, -5116, 6162, 5666, -5657, -6171, 5107, 6624, -4519, -7026, 3896, 7370, -3246, -7657, 2569, 7882, -1877, -8048, 1170, 8150, -457, -8191, -259, 8167, 970, -8084, -1673, 7938, 2361, -7734, -3030, 7472, 3674, -7156, -4291, 6786, 4873, -6369, -5419, 5905, 5923, -5400, -6384, 4856, 6796, -4280, -7160, 3672, 7470, -3042, -7727, 2390, 7928, -1725, -8073, 1047, 8160, -365, -8191, -319, 8164, 998, -8082, -1670, 7943, 2326, -7751, -2968, 7505, 3585, -7211, -4178, 6868, 4740, -6481, -5271, 6049, 5763, -5581, -6218, 5075, 6629, -4539, -6997, 3973, 7317, -3384, -7590, 2773, 7812, -2148, -7985, 1508, 8104, -863, -8174, 212, 8190, 437, -8156, -1083, 8070, 1719, -7935, -2344, 7750, 2951, -7520, -3541, 7242, 4105, -6923, -4645, 6561, 5154, -6162, -5632, 5726, 6073, -5259, -6479, 4759, 6843, -4236, -7169, 3686, 7449, -3119, -7688, 2534, 7879, -1937, -8027, 1329, 8126, -717, -8181, 101, 8188, 512, -8151, -1123, 8066, 1723, -7938, -2315, 7766, 2890, -7553, -3449, 7297, 3986, -7004, -4502, 6673, 4990, -6309, -5452, 5910, 5882, -5482, -6282, 5026, 6645, -4546, -6974, 4042, 7265, -3520, -7518, 2980, 7731, -2428, -7905, 1863, 8037, -1293, -8130, 715, 8179, -138, -8190, -440, 8158, 1012, -8088, -1579, 7977, 2136, -7829, -2682, 7642, 3211, -7420, -3725, 7162, 4219, -6872, -4692, 6549, 5140, -6198, -5565, 5817, 5960, -5413, -6329, 4982, 6665, -4533, -6972, 4062, 7245, -3576, -7486, 3073, 7690, -2561, -7862, 2037, 7996, -1507, -8097, 971, 8160, -434, -8190, -106, 8182, 641, -8141, -1173, 8064, 1697, -7954, -2214, 7810, 2718, -7635, -3211, 7428, 3687, -7192, -4149, 6926, 4590, -6635, -5013, 6315, 5412, -5974, -5791, 5608, 6143, -5222, -6472, 4816, 6772, -4394, -7047, 3954, 7292, -3503, -7510, 3038, 7696, -2565, -7855, 2082, 7982, -1594, -8080, 1101, 8146, -607, -8184, 110, 8189, 383, -8167, -875, 8114, 1360, -8033, -1841, 7923, 2311, -7786, -2774, 7621, 3223, -7432, -3662, 7216, 4084, -6978, -4493, 6715, 4883, -6432, -5257, 6127, 5610, -5804, -5945, 5461, 6258, -5104, -6551, 4729, 6819, -4342, -7066, 3941, 7288, -3531, -7488, 3109, 7662, -2681, -7812, 2244, 7936, -1803, -8038, 1357, 8112, -911, -8163, 461, 8187, -14, -8189, -434, 8164, 876, -8118, -1317, 8046, 1749, -7953, -2177, 7835, 2595, -7697, -3006, 7537, 3405, -7357, -3795, 7156, 4171, -6938, -4535, 6700, 4884, -6446, -5221, 6174, 5539, -5889, -5844, 5587, 6130, -5274, -6401, 4946, 6652, -4609, -6887, 4259, 7101, -3902, -7298, 3535, 7475, -3162, -7633, 2781, 7770, -2397, -7890, 2006, 7988, -1614, -8068, 1218, 8127, -823, -8168, 426, 8187, -32, -8190, -363, 8171, 754, -8136, -1143, 8081, 1525, -8010, -1905, 7919, 2276, -7813, -2643, 7689, 3001, -7550, -3352, 7394, 3693, -7225, -4026, 7039, 4347, -6841, -4660, 6628, 4960, -6405, -5250, 6168, 5526, -5921, -5792, 5661, 6043, -5394, -6283, 5115, 6508, -4830, -6720, 4535, 6918, -4235, -7103, 3926, 7271, -3613, -7428, 3293, 7568, -2971, -7695, 2643, 7807, -2313, -7905, 1980, 7987, -1646, -8057, 1309, 8111, -974, -8152, 637, 8177, -302, -8190, -33, 8188, 364, -8174, -696, 8145, 1022, -8105, -1347, 8051, 1666, -7986, -1983, 7906, 2293, -7817, -2600, 7715, 2899, -7603, -3195, 7479, 3482, -7346, -3764, 7202, 4037, -7049, -4305, 6886, 4563, -6715, -4816, 6535, 5058, -6348, -5294, 6151, 5520, -5950, -5738, 5739, 5946, -5525, -6147, 5302, 6337, -5076, -6519, 4842, 6691, -4606, -6854, 4364, 7007, -4119, -7151, 3869, 7285, -3618, -7410, 3362, 7525, -3106, -7632, 2846, 7727, -2586, -7815, 2323, 7892, -2061, -7961, 1796, 8019, -1534, -8071, 1269, 8111, -1006, -8145, 742, 8168, -481, -8184, 220, 8190, 38, -8190, -297, 8180, 551, -8163, -805, 8137, 1055, -8106, -1304, 8065, 1548, -8019, -1791, 7965, 2028, -7905, -2265, 7837, 2495, -7765, -2724, 7684, 2946, -7600, -3167, 7507, 3381, -7412, -3593, 7309, 3799, -7203, -4002, 7090, 4199, -6975, -4392, 6853, 4579, -6729, -4763, 6598, 4940, -6467, -5115, 6329, 5282, -6190, -5446, 6046, 5603, -5901, -5757, 5752, 5904, -5601, -6048, 5447, 6185, -5292, -6319, 5133, 6446, -4974, -6569, 4812, 6686, -4650, -6800, 4484, 6907, -4320, -7011, 4153, 7108, -3987, -7202, 3818, 7290, -3650, -7375, 3481, 7453, -3313, -7529, 3142, 7598, -2974, -7665, 2804, 7725, -2637, -7784, 2468, 7836, -2301, -7886, 2133, 7930, -1967, -7972, 1801, 8008, -1637, -8043, 1472, 8071, -1311, -8099, 1148, 8120, -989, -8141, 829, 8156, -673, -8170, 516, 8179, -363, -8187, 209, 8189, -59, -8191, -92, 8189, 238, -8186, -385, 8178, 528, -8170, -671, 8157, 810, -8144, -950, 8127, 1085, -8110, -1220, 8089, 1351, -8068, -1482, 8043, 1609, -8019, -1736, 7991, 1859, -7963, -1982, 7932, 2101, -7902, -2219, 7868, 2333, -7835, -2447, 7799, 2557, -7764, -2667, 7726, 2773, -7689, -2879, 7649, 2980, -7610, -3081, 7569, 3178, -7529, -3275, 7487, 3368, -7446, -3461, 7402, 3550, -7361, -3638, 7317, 3723, -7275, -3808, 7230, 3888, -7188, -3969, 7143, 4045, -7101, -4122, 7056, 4194, -7014, -4267, 6970, 4336, -6928, -4405, 6884, 4470, -6843, -4535, 6800, 4596, -6759, -4658, 6717, 4716, -6677, -4774, 6636, 4828, -6597, -4882, 6557, 4933, -6520, -4984, 6481, 5032, -6445, -5080, 6408, 5124, -6373, -5168, 6337, 5209, -6304, -5251, 6270, 5289, -6239, -5327, 6206, 5362, -6177, -5398, 6146, 5430, -6119, -5462, 6090, 5491, -6065, -5521, 6038, 5547, -6015, -5574, 5990, 5598, -5969, -5622, 5946, 5643, -5927, -5664, 5907, 5683, -5890, -5702, 5873, 5717, -5858, -5734, 5843, 5747, -5830, -5761, 5817, 5771, -5807, -5782, 5797, 5791, -5789, -5799, 5781, 5805, -5776, -5811, 5770, 5815, -5768, -5819, 5764, 5819, -5764, -5821, 5763, 5819, -5765, -5818, 5767, 5814, -5772, -5811, 5776, 5804, -5783, -5798, 5789, 5789, -5799, -5781, 5808, 5770, -5820, -5759, 5831, 5745, -5846, -5731, 5859, 5715, -5876, -5699, 5892, 5680, -5911, -5662, 5929, 5640, -5950, -5619, 5971, 5594, -5994, -5571, 6017, 5543, -6043, -5517, 6067, 5487, -6095, -5458, 6122, 5425, -6152, -5393, 6180, 5357, -6212, -5322, 6242, 5283, -6276, -5245, 6308, 5203, -6343, -5162, 6377, 5117, -6414, -5073, 6449, 5025, -6487, -4977, 6524, 4926, -6564, -4875, 6602, 4820, -6643, -4765, 6682, 4707, -6724, -4649, 6764, 4587, -6807, -4526, 6848, 4460, -6891, -4395, 6933, 4326, -6977, -4257, 7019, 4184, -7064, -4111, 7106, 4034, -7151, -3957, 7193, 3877, -7238, -3796, 7280, 3711, -7324, -3626, 7366, 3537, -7409, -3448, 7451, 3355, -7494, -3262, 7534, 3164, -7576, -3067, 7615, 2965, -7655, -2864, 7693, 2758, -7732, -2652, 7768, 2542, -7805, -2431, 7839, 2317, -7874, -2202, 7905, 2083, -7937, -1965, 7966, 1842, -7996, -1718, 8022, 1591, -8048, -1464, 8070, 1332, -8093, -1201, 8112, 1065, -8130, -930, 8145, 790, -8160, -651, 8170, 507, -8180, -364, 8185, 217, -8190, -70, 8190, -81, -8190, 231, 8185, -385, -8178, 539, 8167, -696, -8155, 852, 8137, -1012, -8118, 1172, 8094, -1334, -8068, 1496, 8037, -1661, -8004, 1825, 7965, -1991, -7925, 2157, 7878, -2325, -7829, 2492, 7775, -2661, -7718, 2829, 7655, -2999, -7589, 3167, 7517, -3337, -7443, 3505, 7362, -3675, -7278, 3842, 7188, -4011, -7095, 4177, 6995, -4344, -6893, 4508, 6783, -4673, -6671, 4835, 6551, -4997, -6429, 5156, 6299, -5314, -6167, 5469, 6027, -5623, -5884, 5773, 5735, -5923, -5582, 6067, 5422, -6211, -5259, 6349, 5089, -6486, -4916, 6617, 4736, -6747, -4553, 6870, 4364, -6992, -4171, 7106, 3972, -7219, -3770, 7324, 3562, -7426, -3352, 7521, 3135, -7612, -2915, 7696, 2690, -7776, -2463, 7847, 2230, -7914, -1995, 7973, 1755, -8027, -1514, 8072, 1267, -8111, -1020, 8142, 768, -8166, -516, 8181, 259, -8190, -2, 8190, -258, -8182, 518, 8165, -781, -8141, 1043, 8106, -1308, -8064, 1571, 8011, -1836, -7952, 2098, 7881, -2362, -7803, 2623, 7714, -2885, -7617, 3143, 7509, -3400, -7393, 3654, 7266, -3906, -7131, 4154, 6985, -4400, -6831, 4640, 6666, -4877, -6494, 5108, 6310, -5335, -6119, 5555, 5917, -5771, -5708, 5978, 5488, -6181, -5261, 6374, 5024, -6562, -4780, 6740, 4526, -6911, -4267, 7071, 3998, -7224, -3724, 7365, 3440, -7499, -3153, 7619, 2856, -7731, -2556, 7830, 2249, -7919, -1938, 7995, 1620, -8060, -1300, 8111, 975, -8151, -648, 8176, 316, -8190, 15, 8188, -351, -8175, 686, 8146, -1023, -8105, 1358, 8047, -1695, -7977, 2028, 7891, -2361, -7792, 2690, 7677, -3018, -7549, 3339, 7405, -3659, -7249, 3970, 7076, -4278, -6891, 4578, 6690, -4872, -6477, 5156, 6248, -5433, -6008, 5699, 5753, -5957, -5488, 6202, 5208, -6438, -4918, 6660, 4615, -6871, -4302, 7066, 3978, -7250, -3645, 7417, 3301, -7571, -2951, 7707, 2590, -7830, -2224, 7933, 1849, -8021, -1471, 8090, 1086, -8143, -698, 8175, 306, -8191, 88, 8186, -484, -8163, 880, 8119, -1277, -8058, 1670, 7975, -2064, -7874, 2451, 7752, -2837, -7612, 3215, 7450, -3589, -7271, 3953, 7071, -4311, -6854, 4657, 6617, -4995, -6363, 5319, 6090, -5632, -5801, 5930, 5494, -6215, -5173, 6483, 4835, -6736, -4484, 6970, 4117, -7187, -3740, 7383, 3348, -7562, -2948, 7718, 2535, -7854, -2116, 7967, 1687, -8058, -1253, 8125, 812, -8170, -369, 8189, -79, -8186, 526, 8156, -975, -8103, 1422, 8024, -1867, -7921, 2307, 7791, -2743, -7639, 3170, 7460, -3591, -7259, 4000, 7031, -4399, -6782, 4784, 6509, -5157, -6215, 5512, 5897, -5852, -5561, 6172, 5203, -6474, -4828, 6754, 4434, -7014, -4025, 7249, 3598, -7461, -3160, 7647, 2707, -7808, -2245, 7940, 1771, -8047, -1291, 8123, 803, -8172, -313, 8190, -183, -8180, 677, 8138, -1173, -8068, 1664, 7965, -2153, -7834, 2633, 7671, -3107, -7480, 3568, 7258, -4020, -7009, 4455, 6730, -4877, -6426, 5278, 6094, -5663, -5738, 6024, 5356, -6364, -4953, 6678, 4527, -6967, -4084, 7227, 3620, -7461, -3141, 7662, 2646, -7834, -2140, 7971, 1622, -8078, -1097, 8148, 563, -8186, -28, 8187, -511, -8154, 1048, 8084, -1584, -7980, 2113, 7839, -2636, -7664, 3147, 7452, -3647, -7208, 4131, 6929, -4599, -6620, 5046, 6277, -5473, -5906, 5874, 5504, -6250, -5078, 6597, 4624, -6916, -4149, 7201, 3651, -7454, -3136, 7671, 2603, -7853, -2057, 7995, 1497, -8101, -931, 8165, 356, -8191, 221, 8175, -800, -8119, 1375, 8020, -1946, -7883, 2507, 7703, -3059, -7484, 3596, 7225, -4117, -6929, 4616, 6594, -5094, -6226, 5545, 5822, -5970, -5388, 6362, 4921, -6724, -4429, 7048, 3910, -7337, -3370, 7585, 2807, -7794, -2230, 7959, 1637, -8082, -1035, 8158, 424, -8191, 190, 8175, -806, -8116, 1417, 8008, -2024, -7855, 2619, 7655, -3202, -7412, 3767, 7123, -4313, -6794, 4833, 6422, -5328, -6012, 5791, 5564, -6222, -5083, 6615, 4568, -6972, -4026, 7285, 3456, -7556, -2866, 7780, 2254, -7958, -1628, 8085, 989, -8164, -344, 8190, -307, -8167, 956, 8090, -1602, -7963, 2238, 7783, -2863, -7554, 3469, 7273, -4057, -6947, 4617, 6572, -5151, -6155, 5650, 5695, -6115, -5197, 6538, 4661, -6921, -4095, 7256, 3497, -7545, -2876, 7781, 2232, -7967, -1574, 8096, 900, -8172, -221, 8190, -464, -8152, 1145, 8055, -1822, -7903, 2485, 7693, -3135, -7429, 3762, 7110, -4365, -6740, 4937, 6319, -5476, -5854, 5974, 5342, -6432, -4792, 6842, 4203, -7205, -3584, 7513, 2934, -7767, -2263, 7962, 1572, -8100, -868, 8174, 155, -8189, 560, 8139, -1273, -8028, 1977, 7854, -2669, -7619, 3340, 7323, -3989, -6971, 4606, 6561, -5190, -6101, 5732, 5589, -6232, -5033, 6681, 4433, -7080, -3799, 7420, 3130, -7703, -2436, 7922, 1719, -8079, -987, 8167, 244, -8191, 500, 8144, -1245, -8031, 1978, 7849, -2699, -7602, 3397, 7289, -4069, -6914, 4706, 6478, -5307, -5988, 5861, 5442, -6368, -4851, 6819, 4214, -7213, -3541, 7544, 2833, -7810, -2100, 8007, 1346, -8135, -580, 8188, -196, -8171, 969, 8078, -1737, -7914, 2489, 7676, -3222, -7369, 3925, 6992, -4596, -6552, 5224, 6049, -5807, -5491, 6336, 4878, -6808, -4221, 7216, 3520, -7559, -2786, 7829, 2023, -8027, -1241, 8147, 443, -8191, 359, 8155, -1161, -8042, 1952, 7849, -2727, -7580, 3475, 7235, -4193, -6821, 4869, 6336, -5500, -5789, 6077, 5181, -6595, -4523, 7047, 3815, -7431, -3070, 7738, 2290, -7970, -1487, 8119, 666, -8188, 163, 8170, -993, -8070, 1813, 7885, -2617, -7619, 3394, 7271, -4139, -6848, 4840, 6350, -5494, -5786, 6089, 5157, -6622, -4474, 7083, 3740, -7472, -2966, 7778, 2157, -8004, -1324, 8141, 474, -8191, 381, 8150, -1236, -8022, 2077, 7802, -2899, -7498, 3688, 7108, -4440, -6640, 5141, 6094, -5788, -5481, 6370, 4803, -6882, -4070, 7315, 3288, -7667, -2469, 7931, 1618, -8105, -749, 8185, -133, -8171, 1013, 8061, -1885, -7858, 2734, 7561, -3555, -7176, 4334, 6703, -5065, -6153, 5735, 5525, -6340, -4833, 6868, 4079, -7317, -3277, 7676, 2431, -7944, -1556, 8115, 659, -8189, 246, 8161, -1152, -8034, 2043, 7805, -2913, -7482, 3746, 7063, -4536, -6557, 5269, 5965, -5939, -5300, 6533, 4564, -7048, -3771, 7472, 2926, -7804, -2045, 8034, 1134, -8164, -208, 8186, -724, -8105, 1646, 7916, -2551, -7626, 3422, 7233, -4251, -6747, 5025, 6168, -5735, -5509, 6369, 4774, -6921, -3976, 7379, 3121, -7742, -2224, 7999, 1294, -8150, -347, 8189, -608, -8120, 1555, 7937, -2485, -7647, 3380, 7249, -4232, -6753, 5025, 6160, -5752, -5483, 6398, 4726, -6958, -3904, 7419, 3023, -7779, -2100, 8028, 1144, -8165, -171, 8184, -807, -8089, 1773, 7876, -2718, -7551, 3623, 7114, -4480, -6576, 5271, 5940, -5989, -5217, 6618, 4416, -7154, -3550, 7583, 2628, -7904, -1668, 8106, 679, -8190, 319, 8149, -1317, -7989, 2294, 7707, -3240, -7310, 4138, 6800, -4976, -6188, 5738, 5479, -6416, -4687, 6994, 3820, -7469, -2895, 7827, 1921, -8067, -918, 8180, -103, -8169, 1122, 8027, -2127, -7762, 3099, 7372, -4025, -6868, 4887, 6252, -5676, -5537, 6373, 4732, -6972, -3851, 7458, 2905, -7828, -1913, 8069, 886, -8183, 154, 8163, -1196, -8011, 2218, 7726, -3208, -7317, 4144, 6784, -5016, -6141, 5805, 5393, -6500, -4556, 7087, 3640, -7558, -2664, 7902, 1639, -8115, -588, 8190, -478, -8129, 1535, 7928, -2569, -7594, 3560, 7128, -4493, -6541, 5349, 5839, -6116, -5037, 6776, 4144, -7323, -3181, 7741, 2158, -8027, -1099, 8171, 16, -8175, 1067, 8032, -2134, -7749, 3164, 7327, -4141, -6776, 5044, 6102, -5860, -5319, 6571, 4438, -7167, -3478, 7633, 2451, -7963, -1380, 8148, 281, -8187, 823, 8075, -1916, -7817, 2973, 7413, -3979, -6873, 4912, 6205, -5757, -5422, 6495, 4535, -7115, -3565, 7601, 2524, -7947, -1436, 8143, 318, -8188, 806, 8076, -1919, -7813, 2995, 7398, -4017, -6845, 4962, 6157, -5816, -5352, 6557, 4441, -7175, -3445, 7653, 2379, -7985, -1266, 8161, 126, -8179, 1017, 8036, -2143, -7737, 3227, 7283, -4251, -6686, 5191, 5954, -6031, -5105, 6750, 4151, -7337, -3114, 7777, 2012, -8063, -869, 8185, -295, -8145, 1452, 7937, -2584, -7569, 3663, 7045, -4671, -6378, 5582, 5578, -6383, -4664, 7051, 3650, -7577, -2561, 7944, 1416, -8149, -241, 8183, -942, -8048, 2105, 7742, -3228, -7275, 4282, 6652, -5250, -5890, 6106, 4999, -6836, -4004, 7419, 2919, -7846, -1773, 8105, 584, -8191, 616, 8100, -1807, -7835, 2958, 7399, -4049, -6803, 5052, 6056, -5948, -5178, 6712, 4183, -7333, -3097, 7792, 1939, -8081, -739, 8189, -482, -8119, 1691, 7865, -2866, -7438, 3977, 6842, -5003, -6093, 5915, 5205, -6698, -4199, 7328, 3096, -7795, -1922, 8084, 701, -8191, 535, 8109, -1763, -7843, 2951, 7395, -4074, -6777, 5102, 6000, -6016, -5085, 6790, 4049, -7409, -2919, 7854, 1717, -8117, -475, 8189, -781, -8070, 2019, 7759, -3213, -7266, 4330, 6598, -5348, -5774, 6238, 4809, -6983, -3730, 7559, 2558, -7957, -1325, 8161, 57, -8171, 1213, 7981, -2457, -7599, 3641, 7030, -4739, -6291, 5722, 5394, -6568, -4366, 7251, 3228, -7759, -2010, 8074, 739, -8191, 550, 8103, -1829, -7815, 3063, 7330, -4223, -6663, 5277, 5826, -6202, -4843, 6970, 3734, -7564, -2532, 7966, 1262, -8169, 40, 8161, -1345, -7947, 2615, 7528, -3821, -6916, 4929, 6124, -5914, -5175, 6744, 4089, -7404, -2897, 7870, 1627, -8133, -314, 8183, -1010, -8021, 2308, 7646, -3549, -7071, 4695, 6307, -5722, -5377, 6596, 4302, -7298, -3113, 7805, 1837, -8106, -513, 8189, -829, -8054, 2148, 7701, -3413, -7141, 4586, 6386, -5638, -5458)        
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L32_i
    );

    L32C31_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (2123, 8056, -820, -8190, -505, 8107, 1814, -7816, -3075, 7319, 4253, -6636, -5321, 5779, 6249, -4777, -7016, 3651, 7600, -2435, -7991, 1157, 8175, 148, -8152, -1449, 7920, 2710, -7490, -3902, 6869, 4992, -6077, -5957, 5132, 6769, -4061, -7413, 2888, 7868, -1647, -8129, 364, 8186, 924, -8041, -2190, 7696, 3398, -7164, -4522, 6454, 5532, -5589, -6408, 4586, 7123, -3475, -7666, 2279, 8021, -1031, -8182, -242, 8143, 1505, -7911, -2733, 7486, 3891, -6885, -4957, 6118, 5901, -5209, -6705, 4174, 7347, -3044, -7816, 1842, 8098, -600, -8191, -656, 8090, 1894, -7801, -3087, 7329, 4205, -6688, -5225, 5892, 6121, -4961, -6876, 3916, 7470, -2784, -7893, 1587, 8132, -358, -8187, -880, 8054, 2094, -7739, -3261, 7247, 4350, -6594, -5342, 5791, 6210, -4861, -6939, 3822, 7510, -2700, -7914, 1518, 8139, -305, -8186, -914, 8049, 2109, -7737, -3259, 7252, 4333, -6611, -5312, 5825, 6172, -4914, -6899, 3896, 7472, -2796, -7884, 1636, 8124, -444, -8190, -758, 8078, 1940, -7795, -3081, 7344, 4152, -6739, -5136, 5990, 6007, -5117, -6752, 4135, 7351, -3069, -7797, 1939, 8077, -772, -8190, -412, 8129, 1584, -7902, -2722, 7509, 3801, -6964, -4802, 6274, 5701, -5458, -6483, 4530, 7130, -3512, -7632, 2422, 7977, -1287, -8161, 125, 8178, 1035, -8032, -2175, 7723, 3267, -7261, -4295, 6654, 5233, -5916, -6068, 5061, 6780, -4108, -7358, 3074, 7789, -1983, -8067, 852, 8186, 291, -8146, -1429, 7946, 2536, -7593, -3594, 7093, 4578, -6458, -5475, 5698, 6264, -4832, -6933, 3873, 7467, -2843, -7860, 1759, 8101, -645, -8191, -481, 8124, 1595, -7907, -2678, 7539, 3708, -7033, -4670, 6395, 5541, -5641, -6310, 4782, 6959, -3838, -7480, 2823, 7862, -1760, -8101, 664, 8190, 441, -8131, -1537, 7923, 2602, -7574, -3621, 7088, 4570, -6476, -5439, 5747, 6206, -4919, -6864, 4003, 7396, -3019, -7799, 1981, 8061, -912, -8183, -174, 8159, 1252, -7995, -2310, 7689, 3323, -7252, -4279, 6688, 5157, -6011, -5947, 5230, 6632, -4363, -7204, 3420, 7650, -2422, -7967, 1383, 8146, -324, -8189, -741, 8092, 1789, -7861, -2808, 7497, 3776, -7010, -4682, 6405, 5506, -5697, -6240, 4894, 6868, -4014, -7383, 3067, 7775, -2073, -8041, 1046, 8174, -5, -8175, -1037, 8042, 2058, -7782, -3046, 7395, 3982, -6892, -4854, 6278, 5645, -5567, -6348, 4767, 6947, -3895, -7437, 2961, 7807, -1984, -8056, 975, 8177, 45, -8173, -1064, 8039, 2064, -7784, -3032, 7406, 3949, -6918, -4807, 6323, 5587, -5634, -6283, 4858, 6880, -4012, -7375, 3105, 7755, -2155, -8020, 1173, 8163, -176, -8185, -824, 8084, 1807, -7865, -2765, 7528, 3677, -7083, -4537, 6533, 5326, -5890, -6038, 5161, 6659, -4360, -7185, 3495, 7604, -2584, -7914, 1635, 8109, -666, -8190, -313, 8151, 1283, -8000, -2236, 7733, 3153, -7360, -4026, 6882, 4840, -6311, -5586, 5651, 6251, -4916, -6831, 4111, 7313, -3254, -7695, 2352, 7970, -1420, -8137, 470, 8190, 484, -8135, -1431, 7968, 2355, -7696, -3248, 7319, 4094, -6846, -4885, 6282, 5609, -5637, -6258, 4917, 6822, -4135, -7297, 3298, 7673, -2422, -7951, 1514, 8122, -590, -8191, -342, 8151, 1266, -8008, -2174, 7761, 3051, -7418, -3889, 6978, 4674, -6453, -5400, 5846, 6055, -5168, -6635, 4425, 7129, -3629, -7535, 2789, 7844, -1917, -8058, 1021, 8171, -116, -8185, -790, 8096, 1683, -7912, -2556, 7629, 3394, -7257, -4192, 6796, 4936, -6257, -5621, 5642, 6236, -4963, -6778, 4224, 7236, -3439, -7610, 2613, 7892, -1760, -8084, 886, 8178, -6, -8180, -875, 8085, 1742, -7899, -2590, 7621, 3404, -7258, -4179, 6812, 4904, -6291, -5574, 5698, 6177, -5044, -6712, 4333, 7169, -3577, -7548, 2781, 7839, -1958, -8046, 1112, 8162, -259, -8190, -598, 8126, 1445, -7977, -2276, 7739, 3079, -7420, -3850, 7021, 4575, -6549, -5252, 6006, 5870, -5403, -6427, 4742, 6912, -4034, -7327, 3284, 7661, -2502, -7917, 1695, 8089, -873, -8179, 43, 8182, 785, -8104, -1605, 7941, 2404, -7700, -3180, 7379, 3920, -6987, -4621, 6523, 5272, -5998, -5872, 5412, 6409, -4775, -6885, 4091, 7290, -3370, -7624, 2615, 7881, -1839, -8063, 1045, 8165, -244, -8190, -559, 8134, 1354, -8003, -2136, 7794, 2893, -7514, -3624, 7161, 4317, -6744, -4971, 6263, 5574, -5726, -6126, 5136, 6619, -4502, -7052, 3826, 7417, -3118, -7715, 2381, 7941, -1627, -8097, 857, 8177, -84, -8186, -691, 8120, 1456, -7984, -2208, 7775, 2937, -7501, -3640, 7159, 4308, -6758, -4939, 6297, 5524, -5785, -6062, 5222, 6545, -4617, -6972, 3973, 7338, -3298, -7642, 2595, 7879, -1874, -8052, 1137, 8155, -394, -8191, -353, 8158, 1093, -8060, -1824, 7894, 2537, -7666, -3229, 7374, 3892, -7026, -4523, 6619, 5115, -6163, -5667, 5656, 6170, -5108, -6625, 4518, 7025, -3897, -7371, 3245, 7656, -2570, -7883, 1876, 8047, -1171, -8151, 456, 8190, 258, -8168, -971, 8083, 1672, -7939, -2362, 7733, 3029, -7473, -3675, 7155, 4290, -6787, -4874, 6368, 5418, -5906, -5924, 5399, 6383, -4857, -6797, 4279, 7159, -3673, -7471, 3041, 7726, -2391, -7929, 1724, 8072, -1048, -8161, 364, 8190, 318, -8165, -999, 8081, 1669, -7944, -2327, 7750, 2967, -7506, -3586, 7210, 4177, -6869, -4741, 6480, 5270, -6050, -5764, 5580, 6217, -5076, -6630, 4538, 6996, -3974, -7318, 3383, 7589, -2774, -7813, 2147, 7984, -1509, -8105, 862, 8173, -213, -8191, -438, 8155, 1082, -8071, -1720, 7934, 2343, -7751, -2952, 7519, 3540, -7243, -4106, 6922, 4644, -6562, -5155, 6161, 5631, -5727, -6074, 5258, 6478, -4760, -6844, 4235, 7168, -3687, -7450, 3118, 7687, -2535, -7880, 1936, 8026, -1330, -8127, 716, 8180, -102, -8189, -513, 8150, 1122, -8067, -1724, 7937, 2314, -7767, -2891, 7552, 3448, -7298, -3987, 7003, 4501, -6674, -4991, 6308, 5451, -5911, -5883, 5481, 6281, -5027, -6646, 4545, 6973, -4043, -7266, 3519, 7517, -2981, -7732, 2427, 7904, -1864, -8038, 1292, 8129, -716, -8180, 137, 8189, 439, -8159, -1013, 8087, 1578, -7978, -2137, 7828, 2681, -7643, -3212, 7419, 3724, -7163, -4220, 6871, 4691, -6550, -5141, 6197, 5564, -5818, -5961, 5412, 6328, -4983, -6666, 4532, 6971, -4063, -7246, 3575, 7485, -3074, -7691, 2560, 7861, -2038, -7997, 1506, 8096, -972, -8161, 433, 8189, 105, -8183, -642, 8140, 1172, -8065, -1698, 7953, 2213, -7811, -2719, 7634, 3210, -7429, -3688, 7191, 4148, -6927, -4591, 6634, 5012, -6316, -5413, 5973, 5790, -5609, -6144, 5221, 6471, -4817, -6773, 4393, 7046, -3955, -7293, 3502, 7509, -3039, -7697, 2564, 7854, -2083, -7983, 1593, 8079, -1102, -8147, 606, 8183, -111, -8190, -384, 8166, 874, -8115, -1361, 8032, 1840, -7924, -2312, 7785, 2773, -7622, -3224, 7431, 3661, -7217, -4085, 6977, 4492, -6716, -4884, 6431, 5256, -6128, -5611, 5803, 5944, -5462, -6259, 5103, 6550, -4730, -6820, 4341, 7065, -3942, -7289, 3530, 7487, -3110, -7663, 2680, 7811, -2245, -7937, 1802, 8037, -1358, -8113, 910, 8162, -462, -8188, 13, 8188, 433, -8165, -877, 8117, 1316, -8047, -1750, 7952, 2176, -7836, -2596, 7696, 3005, -7538, -3406, 7356, 3794, -7157, -4172, 6937, 4534, -6701, -4885, 6445, 5220, -6175, -5540, 5888, 5843, -5588, -6131, 5273, 6400, -4947, -6653, 4608, 6886, -4260, -7102, 3901, 7297, -3536, -7476, 3161, 7632, -2782, -7771, 2396, 7889, -2007, -7989, 1613, 8067, -1219, -8128, 822, 8167, -427, -8188, 31, 8189, 362, -8172, -755, 8135, 1142, -8082, -1526, 8009, 1904, -7920, -2277, 7812, 2642, -7690, -3002, 7549, 3351, -7395, -3694, 7224, 4025, -7040, -4348, 6840, 4659, -6629, -4961, 6404, 5249, -6169, -5527, 5920, 5791, -5662, -6044, 5393, 6282, -5116, -6509, 4829, 6719, -4536, -6919, 4234, 7102, -3927, -7272, 3612, 7427, -3294, -7569, 2970, 7694, -2644, -7808, 2312, 7904, -1981, -7988, 1645, 8056, -1310, -8112, 973, 8151, -638, -8178, 301, 8189, 32, -8189, -365, 8173, 695, -8146, -1023, 8104, 1346, -8052, -1667, 7985, 1982, -7907, -2294, 7816, 2599, -7716, -2900, 7602, 3194, -7480, -3483, 7345, 3763, -7203, -4038, 7048, 4304, -6887, -4564, 6714, 4815, -6536, -5059, 6347, 5293, -6152, -5521, 5949, 5737, -5740, -5947, 5524, 6146, -5303, -6338, 5075, 6518, -4843, -6692, 4605, 6853, -4365, -7008, 4118, 7150, -3870, -7286, 3617, 7409, -3363, -7526, 3105, 7631, -2847, -7728, 2585, 7814, -2324, -7893, 2060, 7960, -1797, -8020, 1533, 8070, -1270, -8112, 1005, 8144, -743, -8169, 480, 8183, -221, -8191, -39, 8189, 296, -8181, -552, 8162, 804, -8138, -1056, 8105, 1303, -8066, -1549, 8018, 1790, -7966, -2029, 7904, 2264, -7838, -2496, 7764, 2723, -7685, -2947, 7599, 3166, -7508, -3382, 7411, 3592, -7310, -3800, 7202, 4001, -7091, -4200, 6974, 4391, -6854, -4580, 6728, 4762, -6599, -4941, 6466, 5114, -6330, -5283, 6189, 5445, -6047, -5604, 5900, 5756, -5753, -5905, 5600, 6047, -5448, -6186, 5291, 6318, -5134, -6447, 4973, 6568, -4813, -6687, 4649, 6799, -4485, -6908, 4319, 7010, -4154, -7109, 3986, 7201, -3819, -7291, 3649, 7374, -3482, -7454, 3312, 7528, -3143, -7599, 2973, 7664, -2805, -7726, 2636, 7783, -2469, -7837, 2300, 7885, -2134, -7931, 1966, 7971, -1802, -8009, 1636, 8042, -1473, -8072, 1310, 8098, -1149, -8121, 988, 8140, -830, -8157, 672, 8169, -517, -8180, 362, 8186, -210, -8190, 58, 8190, 91, -8190, -239, 8185, 384, -8179, -529, 8169, 670, -8158, -811, 8143, 949, -8128, -1086, 8109, 1219, -8090, -1352, 8067, 1481, -8044, -1610, 8018, 1735, -7992, -1860, 7962, 1981, -7933, -2102, 7901, 2218, -7869, -2334, 7834, 2446, -7800, -2558, 7763, 2666, -7727, -2774, 7688, 2878, -7650, -2981, 7609, 3080, -7570, -3179, 7528, 3274, -7488, -3369, 7445, 3460, -7403, -3551, 7360, 3637, -7318, -3724, 7274, 3807, -7231, -3889, 7187, 3968, -7144, -4046, 7100, 4121, -7057, -4195, 7013, 4266, -6971, -4337, 6927, 4404, -6885, -4471, 6842, 4534, -6801, -4597, 6758, 4657, -6718, -4717, 6676, 4773, -6637, -4829, 6596, 4881, -6558, -4934, 6519, 4983, -6482, -5033, 6444, 5079, -6409, -5125, 6372, 5167, -6338, -5210, 6303, 5250, -6271, -5290, 6238, 5326, -6207, -5363, 6176, 5397, -6147, -5431, 6118, 5461, -6091, -5492, 6064, 5520, -6039, -5548, 6014, 5573, -5991, -5599, 5968, 5621, -5947, -5644, 5926, 5663, -5908, -5684, 5889, 5701, -5874, -5718, 5857, 5733, -5844, -5748, 5829, 5760, -5818, -5772, 5806, 5781, -5798, -5792, 5788, 5798, -5782, -5806, 5775, 5810, -5771, -5816, 5767, 5818, -5765, -5820, 5763, 5820, -5764, -5820, 5764, 5817, -5768, -5815, 5771, 5810, -5777, -5805, 5782, 5797, -5790, -5790, 5798, 5780, -5809, -5771, 5819, 5758, -5832, -5746, 5845, 5730, -5860, -5716, 5875, 5698, -5893, -5681, 5910, 5661, -5930, -5641, 5949, 5618, -5972, -5595, 5993, 5570, -6018, -5544, 6042, 5516, -6068, -5488, 6094, 5457, -6123, -5426, 6151, 5392, -6181, -5358, 6211, 5321, -6243, -5284, 6275, 5244, -6309, -5204, 6342, 5161, -6378, -5118, 6413, 5072, -6450, -5026, 6486, 4976, -6525, -4927, 6563, 4874, -6603, -4821, 6642, 4764, -6683, -4708, 6723, 4648, -6765, -4588, 6806, 4525, -6849, -4461, 6890, 4394, -6934, -4327, 6976, 4256, -7020, -4185, 7063, 4110, -7107, -4035, 7150, 3956, -7194, -3878, 7237, 3795, -7281, -3712, 7323, 3625, -7367, -3538, 7408, 3447, -7452, -3356, 7493, 3261, -7535, -3165, 7575, 3066, -7616, -2966, 7654, 2863, -7694, -2759, 7731, 2651, -7769, -2543, 7804, 2430, -7840, -2318, 7873, 2201, -7906, -2084, 7936, 1964, -7967, -1843, 7995, 1717, -8023, -1592, 8047, 1463, -8071, -1333, 8092, 1200, -8113, -1066, 8129, 929, -8146, -791, 8159, 650, -8171, -508, 8179, 363, -8186, -218, 8189, 69, -8191, 80, 8189, -232, -8186, 384, 8177, -540, -8168, 695, 8154, -853, -8138, 1011, 8117, -1173, -8095, 1333, 8067, -1497, -8038, 1660, 8003, -1826, -7966, 1990, 7924, -2158, -7879, 2324, 7828, -2493, -7776, 2660, 7717, -2830, -7656, 2998, 7588, -3168, -7518, 3336, 7442, -3506, -7363, 3674, 7277, -3843, -7189, 4010, 7094, -4178, -6996, 4343, 6892, -4509, -6784, 4672, 6670, -4836, -6552, 4996, 6428, -5157, -6300, 5313, 6166, -5470, -6028, 5622, 5883, -5774, -5736, 5922, 5581, -6068, -5423, 6210, 5258, -6350, -5090, 6485, 4915, -6618, -4737, 6746, 4552, -6871, -4365, 6991, 4170, -7107, -3973, 7218, 3769, -7325, -3563, 7425, 3351, -7522, -3136, 7611, 2914, -7697, -2691, 7775, 2462, -7848, -2231, 7913, 1994, -7974, -1756, 8026, 1513, -8073, -1268, 8110, 1019, -8143, -769, 8165, 515, -8182, -260, 8189, 1, -8191, 257, 8181, -519, -8166, 780, 8140, -1044, -8107, 1307, 8063, -1572, -8012, 1835, 7951, -2099, -7882, 2361, 7802, -2624, -7715, 2884, 7616, -3144, -7510, 3399, 7392, -3655, -7267, 3905, 7130, -4155, -6986, 4399, 6830, -4641, -6667, 4876, 6493, -5109, -6311, 5334, 6118, -5556, -5918, 5770, 5707, -5979, -5489, 6180, 5260, -6375, -5025, 6561, 4779, -6741, -4527, 6910, 4266, -7072, -3999, 7223, 3723, -7366, -3441, 7498, 3152, -7620, -2857, 7730, 2555, -7831, -2250, 7918, 1937, -7996, -1621, 8059, 1299, -8112, -976, 8150, 647, -8177, -317, 8189, -16, -8189, 350, 8174, -687, -8147, 1022, 8104, -1359, -8048, 1694, 7976, -2029, -7892, 2360, 7791, -2691, -7678, 3017, 7548, -3340, -7406, 3658, 7248, -3971, -7077, 4277, 6890, -4579, -6691, 4871, 6476, -5157, -6249, 5432, 6007, -5700, -5754, 5956, 5487, -6203, -5209, 6437, 4917, -6661, -4616, 6870, 4301, -7067, -3979, 7249, 3644, -7418, -3302, 7570, 2950, -7708, -2591, 7829, 2223, -7934, -1850, 8020, 1470, -8091, -1087, 8142, 697, -8176, -307, 8190, -89, -8187, 483, 8162, -881, -8120, 1276, 8057, -1671, -7976, 2063, 7873, -2452, -7753, 2836, 7611, -3216, -7451, 3588, 7270, -3954, -7072, 4310, 6853, -4658, -6618, 4994, 6362, -5320, -6091, 5631, 5800, -5931, -5495, 6214, 5172, -6484, -4836, 6735, 4483, -6971, -4118, 7186, 3739, -7384, -3349, 7561, 2947, -7719, -2536, 7853, 2115, -7968, -1688, 8057, 1252, -8126, -813, 8169, 368, -8190, 78, 8185, -527, -8157, 974, 8102, -1423, -8025, 1866, 7920, -2308, -7792, 2742, 7638, -3171, -7461, 3590, 7258, -4001, -7032, 4398, 6781, -4785, -6510, 5156, 6214, -5513, -5898, 5851, 5560, -6173, -5204, 6473, 4827, -6755, -4435, 7013, 4024, -7250, -3599, 7460, 3159, -7648, -2708, 7807, 2244, -7941, -1772, 8046, 1290, -8124, -804, 8171, 312, -8191, 182, 8179, -678, -8139, 1172, 8067, -1665, -7966, 2152, 7833, -2634, -7672, 3106, 7479, -3569, -7259, 4019, 7008, -4456, -6731, 4876, 6425, -5279, -6095, 5662, 5737, -6025, -5357, 6363, 4952, -6679, -4528, 6966, 4083, -7228, -3621, 7460, 3140, -7663, -2647, 7833, 2139, -7972, -1623, 8077, 1096, -8149, -564, 8185, 27, -8188, 510, 8153, -1049, -8085, 1583, 7979, -2114, -7840, 2635, 7663, -3148, -7453, 3646, 7207, -4132, -6930, 4598, 6619, -5047, -6278, 5472, 5905, -5875, -5505, 6249, 5077, -6598, -4625, 6915, 4148, -7202, -3652, 7453, 3135, -7672, -2604, 7852, 2056, -7996, -1498, 8100, 930, -8166, -357, 8190, -222, -8176, 799, 8118, -1376, -8021, 1945, 7882, -2508, -7704, 3058, 7483, -3597, -7226, 4116, 6928, -4617, -6595, 5093, 6225, -5546, -5823, 5969, 5387, -6363, -4922, 6723, 4428, -7049, -3911, 7336, 3369, -7586, -2808, 7793, 2229, -7960, -1638, 8081, 1034, -8159, -425, 8190, -191, -8176, 805, 8115, -1418, -8009, 2023, 7854, -2620, -7656, 3201, 7411, -3768, -7124, 4312, 6793, -4834, -6423, 5327, 6011, -5792, -5565, 6221, 5082, -6616, -4569, 6971, 4025, -7286, -3457, 7555, 2865, -7781, -2255, 7957, 1627, -8086, -990, 8163, 343, -8191, 306, 8166, -957, -8091, 1601, 7962, -2239, -7784, 2862, 7553, -3470, -7274, 4056, 6946, -4618, -6573, 5150, 6154, -5651, -5696, 6114, 5196, -6539, -4662, 6920, 4094, -7257, -3498, 7544, 2875, -7782, -2233, 7966, 1573, -8097, -901, 8171, 220, -8191, 463, 8151, -1146, -8056, 1821, 7902, -2486, -7694, 3134, 7428, -3763, -7111, 4364, 6739, -4938, -6320, 5475, 5853, -5975, -5343, 6431, 4791, -6843, -4204, 7204, 3583, -7514, -2935, 7766, 2262, -7963, -1573, 8099, 867, -8175, -156, 8188, -561, -8140, 1272, 8027, -1978, -7855, 2668, 7618, -3341, -7324, 3988, 6970, -4607, -6562, 5189, 6100, -5733, -5590, 6231, 5032, -6682, -4434, 7079, 3798, -7421, -3131, 7702, 2435, -7923, -1720, 8078, 986, -8168, -245, 8190, -501, -8145, 1244, 8030, -1979, -7850, 2698, 7601, -3398, -7290, 4068, 6913, -4707, -6479, 5306, 5987, -5862, -5443, 6367, 4850, -6820, -4215, 7212, 3540, -7545, -2834, 7809, 2099, -8008, -1347, 8134, 579, -8189, 195, 8170, -970, -8079, 1736, 7913, -2490, -7677, 3221, 7368, -3926, -6993, 4595, 6551, -5225, -6050, 5806, 5490, -6337, -4879, 6807, 4220, -7217, -3521, 7558, 2785, -7830, -2024, 8026, 1240, -8148, -444, 8190, -360, -8156, 1160, 8041, -1953, -7850, 2726, 7579, -3476, -7236, 4192, 6820, -4870, -6337, 5499, 5788, -6078, -5182, 6594, 4522, -7048, -3816, 7430, 3069, -7739, -2291, 7969, 1486, -8120, -667, 8187, -164, -8171, 992, 8069, -1814, -7886, 2616, 7618, -3395, -7272, 4138, 6847, -4841, -6351, 5493, 5785, -6090, -5158, 6621, 4473, -7084, -3741, 7471, 2965, -7779, -2158, 8003, 1323, -8142, -475, 8190, -382, -8151, 1235, 8021, -2078, -7803, 2898, 7497, -3689, -7109, 4439, 6639, -5142, -6095, 5787, 5480, -6371, -4804, 6881, 4069, -7316, -3289, 7666, 2468, -7932, -1619, 8104, 748, -8186, 132, 8170, -1014, -8062, 1884, 7857, -2735, -7562, 3554, 7175, -4335, -6704, 5064, 6152, -5736, -5526, 6339, 4832, -6869, -4080, 7316, 3276, -7677, -2432, 7943, 1555, -8116, -660, 8188, -247, -8162, 1151, 8033, -2044, -7806, 2912, 7481, -3747, -7064, 4535, 6556, -5270, -5966, 5938, 5299, -6534, -4565, 7047, 3770, -7473, -2927, 7803, 2044, -8035, -1135, 8163, 207, -8187, 723, 8104, -1647, -7917, 2550, 7625, -3423, -7234, 4250, 6746, -5026, -6169, 5734, 5508, -6370, -4775, 6920, 3975, -7380, -3122, 7741, 2223, -8000, -1295, 8149, 346, -8190, 607, 8119, -1556, -7938, 2484, 7646, -3381, -7250, 4231, 6752, -5026, -6161, 5751, 5482, -6399, -4727, 6957, 3903, -7420, -3024, 7778, 2099, -8029, -1145, 8164, 170, -8185, 806, 8088, -1774, -7877, 2717, 7550, -3624, -7115, 4479, 6575, -5272, -5941, 5988, 5216, -6619, -4417, 7153, 3549, -7584, -2629, 7903, 1667, -8107, -680, 8189, -320, -8150, 1316, 7988, -2295, -7708, 3239, 7309, -4139, -6801, 4975, 6187, -5739, -5480, 6415, 4686, -6995, -3821, 7468, 2894, -7828, -1922, 8066, 917, -8181, 102, 8168, -1123, -8028, 2126, 7761, -3100, -7373, 4024, 6867, -4888, -6253, 5675, 5536, -6374, -4733, 6971, 3850, -7459, -2906, 7827, 1912, -8070, -887, 8182, -155, -8164, 1195, 8010, -2219, -7727, 3207, 7316, -4145, -6785, 5015, 6140, -5806, -5394, 6499, 4555, -7088, -3641, 7557, 2663, -7903, -1640, 8114, 587, -8191, 477, 8128, -1536, -7929, 2568, 7593, -3561, -7129, 4492, 6540, -5350, -5840, 6115, 5036, -6777, -4145, 7322, 3180, -7742, -2159, 8026, 1098, -8172, -17, 8174, -1068, -8033, 2133, 7748, -3165, -7328, 4140, 6775, -5045, -6103, 5859, 5318, -6572, -4439, 7166, 3477, -7634, -2452, 7962, 1379, -8149, -282, 8186, -824, -8076, 1915, 7816, -2974, -7414, 3978, 6872, -4913, -6206, 5756, 5421, -6496, -4536, 7114, 3564, -7602, -2525, 7946, 1435, -8144, -319, 8187, -807, -8077, 1918, 7812, -2996, -7399, 4016, 6844, -4963, -6158, 5815, 5351, -6558, -4442, 7174, 3444, -7654, -2380, 7984, 1265, -8162, -127, 8178, -1018, -8037, 2142, 7736, -3228, -7284, 4250, 6685, -5192, -5955, 6030, 5104, -6751, -4152, 7336, 3113, -7778, -2013, 8062, 868, -8186, 294, 8144, -1453, -7938, 2583, 7568, -3664, -7046, 4670, 6377, -5583, -5579, 6382, 4663, -7052, -3651, 7576, 2560, -7945, -1417, 8148, 240, -8184, 941, 8047, -2106, -7743, 3227, 7274, -4283, -6653, 5249, 5889, -6107, -5000, 6835, 4003, -7420, -2920, 7845, 1772, -8106, -585, 8190, -617, -8101, 1806, 7834, -2959, -7400, 4048, 6802, -5053, -6057, 5947, 5177, -6713, -4184, 7332, 3096, -7793, -1940, 8080, 738, -8190, 481, 8118, -1692, -7866, 2865, 7437, -3978, -6843, 5002, 6092, -5916, -5206, 6697, 4198, -7329, -3097, 7794, 1921, -8085, -702, 8190, -536, -8110, 1762, 7842, -2952, -7396, 4073, 6776, -5103, -6001, 6015, 5084, -6791, -4050, 7408, 2918, -7855, -1718, 8116, 474, -8190, 780, 8069, -2020, -7760, 3212, 7265, -4331, -6599, 5347, 5773, -6239, -4810, 6982, 3729, -7560, -2559, 7956, 1324, -8162, -58, 8170, -1214, -7982, 2456, 7598, -3642, -7031, 4738, 6290, -5723, -5395, 6567, 4365, -7252, -3229, 7758, 2009, -8075, -740, 8190, -551, -8104, 1828, 7814, -3064, -7331, 4222, 6662, -5278, -5827, 6201, 4842, -6971, -3735, 7563, 2531, -7967, -1263, 8168, -41, -8162, 1344, 7946, -2616, -7529, 3820, 6915, -4930, -6125, 5913, 5174, -6745, -4090, 7403, 2896, -7871, -1628, 8132, 313, -8184, 1009, 8020, -2309, -7647, 3548, 7070, -4696, -6308, 5721, 5376, -6597, -4303, 7297, 3112, -7806, -1838, 8105, 512, -8190, 828, 8053, -2149, -7702, 3412, 7140, -4587, -6387, 5637, 5457)         
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L32C31_i
    );

    L32C32_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-2124, -8057, 819, 8189, 504, -8108, -1815, 7815, 3074, -7320, -4254, 6635, 5320, -5780, -6250, 4776, 7015, -3652, -7601, 2434, 7990, -1158, -8176, -149, 8151, 1448, -7921, -2711, 7489, 3901, -6870, -4993, 6076, 5956, -5133, -6770, 4060, 7412, -2889, -7869, 1646, 8128, -365, -8187, -925, 8040, 2189, -7697, -3399, 7163, 4521, -6455, -5533, 5588, 6407, -4587, -7124, 3474, 7665, -2280, -8022, 1030, 8181, 241, -8144, -1506, 7910, 2732, -7487, -3892, 6884, 4956, -6119, -5902, 5208, 6704, -4175, -7348, 3043, 7815, -1843, -8099, 599, 8190, 655, -8091, -1895, 7800, 3086, -7330, -4206, 6687, 5224, -5893, -6122, 4960, 6875, -3917, -7471, 2783, 7892, -1588, -8133, 357, 8186, 879, -8055, -2095, 7738, 3260, -7248, -4351, 6593, 5341, -5792, -6211, 4860, 6938, -3823, -7511, 2699, 7913, -1519, -8140, 304, 8185, 913, -8050, -2110, 7736, 3258, -7253, -4334, 6610, 5311, -5826, -6173, 4913, 6898, -3897, -7473, 2795, 7883, -1637, -8125, 443, 8189, 757, -8079, -1941, 7794, 3080, -7345, -4153, 6738, 5135, -5991, -6008, 5116, 6751, -4136, -7352, 3068, 7796, -1940, -8078, 771, 8189, 411, -8130, -1585, 7901, 2721, -7510, -3802, 6963, 4801, -6275, -5702, 5457, 6482, -4531, -7131, 3511, 7631, -2423, -7978, 1286, 8160, -126, -8179, -1036, 8031, 2174, -7724, -3268, 7260, 4294, -6655, -5234, 5915, 6067, -5062, -6781, 4107, 7357, -3075, -7790, 1982, 8066, -853, -8187, -292, 8145, 1428, -7947, -2537, 7592, 3593, -7094, -4579, 6457, 5474, -5699, -6265, 4831, 6932, -3874, -7468, 2842, 7859, -1760, -8102, 644, 8190, 480, -8125, -1596, 7906, 2677, -7540, -3709, 7032, 4669, -6396, -5542, 5640, 6309, -4783, -6960, 3837, 7479, -2824, -7863, 1759, 8100, -665, -8191, -442, 8130, 1536, -7924, -2603, 7573, 3620, -7089, -4571, 6475, 5438, -5748, -6207, 4918, 6863, -4004, -7397, 3018, 7798, -1982, -8062, 911, 8182, 173, -8160, -1253, 7994, 2309, -7690, -3324, 7251, 4278, -6689, -5158, 6010, 5946, -5231, -6633, 4362, 7203, -3421, -7651, 2421, 7966, -1384, -8147, 323, 8188, 740, -8093, -1790, 7860, 2807, -7498, -3777, 7009, 4681, -6406, -5507, 5696, 6239, -4895, -6869, 4013, 7382, -3068, -7776, 2072, 8040, -1047, -8175, 4, 8174, 1036, -8043, -2059, 7781, 3045, -7396, -3983, 6891, 4853, -6279, -5646, 5566, 6347, -4768, -6948, 3894, 7436, -2962, -7808, 1983, 8055, -976, -8178, -46, 8172, 1063, -8040, -2065, 7783, 3031, -7407, -3950, 6917, 4806, -6324, -5588, 5633, 6282, -4859, -6881, 4011, 7374, -3106, -7756, 2154, 8019, -1174, -8164, 175, 8184, 823, -8085, -1808, 7864, 2764, -7529, -3678, 7082, 4536, -6534, -5327, 5889, 6037, -5162, -6660, 4359, 7184, -3496, -7605, 2583, 7913, -1636, -8110, 665, 8189, 312, -8152, -1284, 7999, 2235, -7734, -3154, 7359, 4025, -6883, -4841, 6310, 5585, -5652, -6252, 4915, 6830, -4112, -7314, 3253, 7694, -2353, -7971, 1419, 8136, -471, -8191, -485, 8134, 1430, -7969, -2356, 7695, 3247, -7320, -4095, 6845, 4884, -6283, -5610, 5636, 6257, -4918, -6823, 4134, 7296, -3299, -7674, 2421, 7950, -1515, -8123, 589, 8190, 341, -8152, -1267, 8007, 2173, -7762, -3052, 7417, 3888, -6979, -4675, 6452, 5399, -5847, -6056, 5167, 6634, -4426, -7130, 3628, 7534, -2790, -7845, 1916, 8057, -1022, -8172, 115, 8184, 789, -8097, -1684, 7911, 2555, -7630, -3395, 7256, 4191, -6797, -4937, 6256, 5620, -5643, -6237, 4962, 6777, -4225, -7237, 3438, 7609, -2614, -7893, 1759, 8083, -887, -8179, 5, 8179, 874, -8086, -1743, 7898, 2589, -7622, -3405, 7257, 4178, -6813, -4905, 6290, 5573, -5699, -6178, 5043, 6711, -4334, -7170, 3576, 7547, -2782, -7840, 1957, 8045, -1113, -8163, 258, 8189, 597, -8127, -1446, 7976, 2275, -7740, -3080, 7419, 3849, -7022, -4576, 6548, 5251, -6007, -5871, 5402, 6426, -4743, -6913, 4033, 7326, -3285, -7662, 2501, 7916, -1696, -8090, 872, 8178, -44, -8183, -786, 8103, 1604, -7942, -2405, 7699, 3179, -7380, -3921, 6986, 4620, -6524, -5273, 5997, 5871, -5413, -6410, 4774, 6884, -4092, -7291, 3369, 7623, -2616, -7882, 1838, 8062, -1046, -8166, 243, 8189, 558, -8135, -1355, 8002, 2135, -7795, -2894, 7513, 3623, -7162, -4318, 6743, 4970, -6264, -5575, 5725, 6125, -5137, -6620, 4501, 7051, -3827, -7418, 3117, 7714, -2382, -7942, 1626, 8096, -858, -8178, 83, 8185, 690, -8121, -1457, 7983, 2207, -7776, -2938, 7500, 3639, -7160, -4309, 6757, 4938, -6298, -5525, 5784, 6061, -5223, -6546, 4616, 6971, -3974, -7339, 3297, 7641, -2596, -7880, 1873, 8051, -1138, -8156, 393, 8190, 352, -8159, -1094, 8059, 1823, -7895, -2538, 7665, 3228, -7375, -3893, 7025, 4522, -6620, -5116, 6162, 5666, -5657, -6171, 5107, 6624, -4519, -7026, 3896, 7370, -3246, -7657, 2569, 7882, -1877, -8048, 1170, 8150, -457, -8191, -259, 8167, 970, -8084, -1673, 7938, 2361, -7734, -3030, 7472, 3674, -7156, -4291, 6786, 4873, -6369, -5419, 5905, 5923, -5400, -6384, 4856, 6796, -4280, -7160, 3672, 7470, -3042, -7727, 2390, 7928, -1725, -8073, 1047, 8160, -365, -8191, -319, 8164, 998, -8082, -1670, 7943, 2326, -7751, -2968, 7505, 3585, -7211, -4178, 6868, 4740, -6481, -5271, 6049, 5763, -5581, -6218, 5075, 6629, -4539, -6997, 3973, 7317, -3384, -7590, 2773, 7812, -2148, -7985, 1508, 8104, -863, -8174, 212, 8190, 437, -8156, -1083, 8070, 1719, -7935, -2344, 7750, 2951, -7520, -3541, 7242, 4105, -6923, -4645, 6561, 5154, -6162, -5632, 5726, 6073, -5259, -6479, 4759, 6843, -4236, -7169, 3686, 7449, -3119, -7688, 2534, 7879, -1937, -8027, 1329, 8126, -717, -8181, 101, 8188, 512, -8151, -1123, 8066, 1723, -7938, -2315, 7766, 2890, -7553, -3449, 7297, 3986, -7004, -4502, 6673, 4990, -6309, -5452, 5910, 5882, -5482, -6282, 5026, 6645, -4546, -6974, 4042, 7265, -3520, -7518, 2980, 7731, -2428, -7905, 1863, 8037, -1293, -8130, 715, 8179, -138, -8190, -440, 8158, 1012, -8088, -1579, 7977, 2136, -7829, -2682, 7642, 3211, -7420, -3725, 7162, 4219, -6872, -4692, 6549, 5140, -6198, -5565, 5817, 5960, -5413, -6329, 4982, 6665, -4533, -6972, 4062, 7245, -3576, -7486, 3073, 7690, -2561, -7862, 2037, 7996, -1507, -8097, 971, 8160, -434, -8190, -106, 8182, 641, -8141, -1173, 8064, 1697, -7954, -2214, 7810, 2718, -7635, -3211, 7428, 3687, -7192, -4149, 6926, 4590, -6635, -5013, 6315, 5412, -5974, -5791, 5608, 6143, -5222, -6472, 4816, 6772, -4394, -7047, 3954, 7292, -3503, -7510, 3038, 7696, -2565, -7855, 2082, 7982, -1594, -8080, 1101, 8146, -607, -8184, 110, 8189, 383, -8167, -875, 8114, 1360, -8033, -1841, 7923, 2311, -7786, -2774, 7621, 3223, -7432, -3662, 7216, 4084, -6978, -4493, 6715, 4883, -6432, -5257, 6127, 5610, -5804, -5945, 5461, 6258, -5104, -6551, 4729, 6819, -4342, -7066, 3941, 7288, -3531, -7488, 3109, 7662, -2681, -7812, 2244, 7936, -1803, -8038, 1357, 8112, -911, -8163, 461, 8187, -14, -8189, -434, 8164, 876, -8118, -1317, 8046, 1749, -7953, -2177, 7835, 2595, -7697, -3006, 7537, 3405, -7357, -3795, 7156, 4171, -6938, -4535, 6700, 4884, -6446, -5221, 6174, 5539, -5889, -5844, 5587, 6130, -5274, -6401, 4946, 6652, -4609, -6887, 4259, 7101, -3902, -7298, 3535, 7475, -3162, -7633, 2781, 7770, -2397, -7890, 2006, 7988, -1614, -8068, 1218, 8127, -823, -8168, 426, 8187, -32, -8190, -363, 8171, 754, -8136, -1143, 8081, 1525, -8010, -1905, 7919, 2276, -7813, -2643, 7689, 3001, -7550, -3352, 7394, 3693, -7225, -4026, 7039, 4347, -6841, -4660, 6628, 4960, -6405, -5250, 6168, 5526, -5921, -5792, 5661, 6043, -5394, -6283, 5115, 6508, -4830, -6720, 4535, 6918, -4235, -7103, 3926, 7271, -3613, -7428, 3293, 7568, -2971, -7695, 2643, 7807, -2313, -7905, 1980, 7987, -1646, -8057, 1309, 8111, -974, -8152, 637, 8177, -302, -8190, -33, 8188, 364, -8174, -696, 8145, 1022, -8105, -1347, 8051, 1666, -7986, -1983, 7906, 2293, -7817, -2600, 7715, 2899, -7603, -3195, 7479, 3482, -7346, -3764, 7202, 4037, -7049, -4305, 6886, 4563, -6715, -4816, 6535, 5058, -6348, -5294, 6151, 5520, -5950, -5738, 5739, 5946, -5525, -6147, 5302, 6337, -5076, -6519, 4842, 6691, -4606, -6854, 4364, 7007, -4119, -7151, 3869, 7285, -3618, -7410, 3362, 7525, -3106, -7632, 2846, 7727, -2586, -7815, 2323, 7892, -2061, -7961, 1796, 8019, -1534, -8071, 1269, 8111, -1006, -8145, 742, 8168, -481, -8184, 220, 8190, 38, -8190, -297, 8180, 551, -8163, -805, 8137, 1055, -8106, -1304, 8065, 1548, -8019, -1791, 7965, 2028, -7905, -2265, 7837, 2495, -7765, -2724, 7684, 2946, -7600, -3167, 7507, 3381, -7412, -3593, 7309, 3799, -7203, -4002, 7090, 4199, -6975, -4392, 6853, 4579, -6729, -4763, 6598, 4940, -6467, -5115, 6329, 5282, -6190, -5446, 6046, 5603, -5901, -5757, 5752, 5904, -5601, -6048, 5447, 6185, -5292, -6319, 5133, 6446, -4974, -6569, 4812, 6686, -4650, -6800, 4484, 6907, -4320, -7011, 4153, 7108, -3987, -7202, 3818, 7290, -3650, -7375, 3481, 7453, -3313, -7529, 3142, 7598, -2974, -7665, 2804, 7725, -2637, -7784, 2468, 7836, -2301, -7886, 2133, 7930, -1967, -7972, 1801, 8008, -1637, -8043, 1472, 8071, -1311, -8099, 1148, 8120, -989, -8141, 829, 8156, -673, -8170, 516, 8179, -363, -8187, 209, 8189, -59, -8191, -92, 8189, 238, -8186, -385, 8178, 528, -8170, -671, 8157, 810, -8144, -950, 8127, 1085, -8110, -1220, 8089, 1351, -8068, -1482, 8043, 1609, -8019, -1736, 7991, 1859, -7963, -1982, 7932, 2101, -7902, -2219, 7868, 2333, -7835, -2447, 7799, 2557, -7764, -2667, 7726, 2773, -7689, -2879, 7649, 2980, -7610, -3081, 7569, 3178, -7529, -3275, 7487, 3368, -7446, -3461, 7402, 3550, -7361, -3638, 7317, 3723, -7275, -3808, 7230, 3888, -7188, -3969, 7143, 4045, -7101, -4122, 7056, 4194, -7014, -4267, 6970, 4336, -6928, -4405, 6884, 4470, -6843, -4535, 6800, 4596, -6759, -4658, 6717, 4716, -6677, -4774, 6636, 4828, -6597, -4882, 6557, 4933, -6520, -4984, 6481, 5032, -6445, -5080, 6408, 5124, -6373, -5168, 6337, 5209, -6304, -5251, 6270, 5289, -6239, -5327, 6206, 5362, -6177, -5398, 6146, 5430, -6119, -5462, 6090, 5491, -6065, -5521, 6038, 5547, -6015, -5574, 5990, 5598, -5969, -5622, 5946, 5643, -5927, -5664, 5907, 5683, -5890, -5702, 5873, 5717, -5858, -5734, 5843, 5747, -5830, -5761, 5817, 5771, -5807, -5782, 5797, 5791, -5789, -5799, 5781, 5805, -5776, -5811, 5770, 5815, -5768, -5819, 5764, 5819, -5764, -5821, 5763, 5819, -5765, -5818, 5767, 5814, -5772, -5811, 5776, 5804, -5783, -5798, 5789, 5789, -5799, -5781, 5808, 5770, -5820, -5759, 5831, 5745, -5846, -5731, 5859, 5715, -5876, -5699, 5892, 5680, -5911, -5662, 5929, 5640, -5950, -5619, 5971, 5594, -5994, -5571, 6017, 5543, -6043, -5517, 6067, 5487, -6095, -5458, 6122, 5425, -6152, -5393, 6180, 5357, -6212, -5322, 6242, 5283, -6276, -5245, 6308, 5203, -6343, -5162, 6377, 5117, -6414, -5073, 6449, 5025, -6487, -4977, 6524, 4926, -6564, -4875, 6602, 4820, -6643, -4765, 6682, 4707, -6724, -4649, 6764, 4587, -6807, -4526, 6848, 4460, -6891, -4395, 6933, 4326, -6977, -4257, 7019, 4184, -7064, -4111, 7106, 4034, -7151, -3957, 7193, 3877, -7238, -3796, 7280, 3711, -7324, -3626, 7366, 3537, -7409, -3448, 7451, 3355, -7494, -3262, 7534, 3164, -7576, -3067, 7615, 2965, -7655, -2864, 7693, 2758, -7732, -2652, 7768, 2542, -7805, -2431, 7839, 2317, -7874, -2202, 7905, 2083, -7937, -1965, 7966, 1842, -7996, -1718, 8022, 1591, -8048, -1464, 8070, 1332, -8093, -1201, 8112, 1065, -8130, -930, 8145, 790, -8160, -651, 8170, 507, -8180, -364, 8185, 217, -8190, -70, 8190, -81, -8190, 231, 8185, -385, -8178, 539, 8167, -696, -8155, 852, 8137, -1012, -8118, 1172, 8094, -1334, -8068, 1496, 8037, -1661, -8004, 1825, 7965, -1991, -7925, 2157, 7878, -2325, -7829, 2492, 7775, -2661, -7718, 2829, 7655, -2999, -7589, 3167, 7517, -3337, -7443, 3505, 7362, -3675, -7278, 3842, 7188, -4011, -7095, 4177, 6995, -4344, -6893, 4508, 6783, -4673, -6671, 4835, 6551, -4997, -6429, 5156, 6299, -5314, -6167, 5469, 6027, -5623, -5884, 5773, 5735, -5923, -5582, 6067, 5422, -6211, -5259, 6349, 5089, -6486, -4916, 6617, 4736, -6747, -4553, 6870, 4364, -6992, -4171, 7106, 3972, -7219, -3770, 7324, 3562, -7426, -3352, 7521, 3135, -7612, -2915, 7696, 2690, -7776, -2463, 7847, 2230, -7914, -1995, 7973, 1755, -8027, -1514, 8072, 1267, -8111, -1020, 8142, 768, -8166, -516, 8181, 259, -8190, -2, 8190, -258, -8182, 518, 8165, -781, -8141, 1043, 8106, -1308, -8064, 1571, 8011, -1836, -7952, 2098, 7881, -2362, -7803, 2623, 7714, -2885, -7617, 3143, 7509, -3400, -7393, 3654, 7266, -3906, -7131, 4154, 6985, -4400, -6831, 4640, 6666, -4877, -6494, 5108, 6310, -5335, -6119, 5555, 5917, -5771, -5708, 5978, 5488, -6181, -5261, 6374, 5024, -6562, -4780, 6740, 4526, -6911, -4267, 7071, 3998, -7224, -3724, 7365, 3440, -7499, -3153, 7619, 2856, -7731, -2556, 7830, 2249, -7919, -1938, 7995, 1620, -8060, -1300, 8111, 975, -8151, -648, 8176, 316, -8190, 15, 8188, -351, -8175, 686, 8146, -1023, -8105, 1358, 8047, -1695, -7977, 2028, 7891, -2361, -7792, 2690, 7677, -3018, -7549, 3339, 7405, -3659, -7249, 3970, 7076, -4278, -6891, 4578, 6690, -4872, -6477, 5156, 6248, -5433, -6008, 5699, 5753, -5957, -5488, 6202, 5208, -6438, -4918, 6660, 4615, -6871, -4302, 7066, 3978, -7250, -3645, 7417, 3301, -7571, -2951, 7707, 2590, -7830, -2224, 7933, 1849, -8021, -1471, 8090, 1086, -8143, -698, 8175, 306, -8191, 88, 8186, -484, -8163, 880, 8119, -1277, -8058, 1670, 7975, -2064, -7874, 2451, 7752, -2837, -7612, 3215, 7450, -3589, -7271, 3953, 7071, -4311, -6854, 4657, 6617, -4995, -6363, 5319, 6090, -5632, -5801, 5930, 5494, -6215, -5173, 6483, 4835, -6736, -4484, 6970, 4117, -7187, -3740, 7383, 3348, -7562, -2948, 7718, 2535, -7854, -2116, 7967, 1687, -8058, -1253, 8125, 812, -8170, -369, 8189, -79, -8186, 526, 8156, -975, -8103, 1422, 8024, -1867, -7921, 2307, 7791, -2743, -7639, 3170, 7460, -3591, -7259, 4000, 7031, -4399, -6782, 4784, 6509, -5157, -6215, 5512, 5897, -5852, -5561, 6172, 5203, -6474, -4828, 6754, 4434, -7014, -4025, 7249, 3598, -7461, -3160, 7647, 2707, -7808, -2245, 7940, 1771, -8047, -1291, 8123, 803, -8172, -313, 8190, -183, -8180, 677, 8138, -1173, -8068, 1664, 7965, -2153, -7834, 2633, 7671, -3107, -7480, 3568, 7258, -4020, -7009, 4455, 6730, -4877, -6426, 5278, 6094, -5663, -5738, 6024, 5356, -6364, -4953, 6678, 4527, -6967, -4084, 7227, 3620, -7461, -3141, 7662, 2646, -7834, -2140, 7971, 1622, -8078, -1097, 8148, 563, -8186, -28, 8187, -511, -8154, 1048, 8084, -1584, -7980, 2113, 7839, -2636, -7664, 3147, 7452, -3647, -7208, 4131, 6929, -4599, -6620, 5046, 6277, -5473, -5906, 5874, 5504, -6250, -5078, 6597, 4624, -6916, -4149, 7201, 3651, -7454, -3136, 7671, 2603, -7853, -2057, 7995, 1497, -8101, -931, 8165, 356, -8191, 221, 8175, -800, -8119, 1375, 8020, -1946, -7883, 2507, 7703, -3059, -7484, 3596, 7225, -4117, -6929, 4616, 6594, -5094, -6226, 5545, 5822, -5970, -5388, 6362, 4921, -6724, -4429, 7048, 3910, -7337, -3370, 7585, 2807, -7794, -2230, 7959, 1637, -8082, -1035, 8158, 424, -8191, 190, 8175, -806, -8116, 1417, 8008, -2024, -7855, 2619, 7655, -3202, -7412, 3767, 7123, -4313, -6794, 4833, 6422, -5328, -6012, 5791, 5564, -6222, -5083, 6615, 4568, -6972, -4026, 7285, 3456, -7556, -2866, 7780, 2254, -7958, -1628, 8085, 989, -8164, -344, 8190, -307, -8167, 956, 8090, -1602, -7963, 2238, 7783, -2863, -7554, 3469, 7273, -4057, -6947, 4617, 6572, -5151, -6155, 5650, 5695, -6115, -5197, 6538, 4661, -6921, -4095, 7256, 3497, -7545, -2876, 7781, 2232, -7967, -1574, 8096, 900, -8172, -221, 8190, -464, -8152, 1145, 8055, -1822, -7903, 2485, 7693, -3135, -7429, 3762, 7110, -4365, -6740, 4937, 6319, -5476, -5854, 5974, 5342, -6432, -4792, 6842, 4203, -7205, -3584, 7513, 2934, -7767, -2263, 7962, 1572, -8100, -868, 8174, 155, -8189, 560, 8139, -1273, -8028, 1977, 7854, -2669, -7619, 3340, 7323, -3989, -6971, 4606, 6561, -5190, -6101, 5732, 5589, -6232, -5033, 6681, 4433, -7080, -3799, 7420, 3130, -7703, -2436, 7922, 1719, -8079, -987, 8167, 244, -8191, 500, 8144, -1245, -8031, 1978, 7849, -2699, -7602, 3397, 7289, -4069, -6914, 4706, 6478, -5307, -5988, 5861, 5442, -6368, -4851, 6819, 4214, -7213, -3541, 7544, 2833, -7810, -2100, 8007, 1346, -8135, -580, 8188, -196, -8171, 969, 8078, -1737, -7914, 2489, 7676, -3222, -7369, 3925, 6992, -4596, -6552, 5224, 6049, -5807, -5491, 6336, 4878, -6808, -4221, 7216, 3520, -7559, -2786, 7829, 2023, -8027, -1241, 8147, 443, -8191, 359, 8155, -1161, -8042, 1952, 7849, -2727, -7580, 3475, 7235, -4193, -6821, 4869, 6336, -5500, -5789, 6077, 5181, -6595, -4523, 7047, 3815, -7431, -3070, 7738, 2290, -7970, -1487, 8119, 666, -8188, 163, 8170, -993, -8070, 1813, 7885, -2617, -7619, 3394, 7271, -4139, -6848, 4840, 6350, -5494, -5786, 6089, 5157, -6622, -4474, 7083, 3740, -7472, -2966, 7778, 2157, -8004, -1324, 8141, 474, -8191, 381, 8150, -1236, -8022, 2077, 7802, -2899, -7498, 3688, 7108, -4440, -6640, 5141, 6094, -5788, -5481, 6370, 4803, -6882, -4070, 7315, 3288, -7667, -2469, 7931, 1618, -8105, -749, 8185, -133, -8171, 1013, 8061, -1885, -7858, 2734, 7561, -3555, -7176, 4334, 6703, -5065, -6153, 5735, 5525, -6340, -4833, 6868, 4079, -7317, -3277, 7676, 2431, -7944, -1556, 8115, 659, -8189, 246, 8161, -1152, -8034, 2043, 7805, -2913, -7482, 3746, 7063, -4536, -6557, 5269, 5965, -5939, -5300, 6533, 4564, -7048, -3771, 7472, 2926, -7804, -2045, 8034, 1134, -8164, -208, 8186, -724, -8105, 1646, 7916, -2551, -7626, 3422, 7233, -4251, -6747, 5025, 6168, -5735, -5509, 6369, 4774, -6921, -3976, 7379, 3121, -7742, -2224, 7999, 1294, -8150, -347, 8189, -608, -8120, 1555, 7937, -2485, -7647, 3380, 7249, -4232, -6753, 5025, 6160, -5752, -5483, 6398, 4726, -6958, -3904, 7419, 3023, -7779, -2100, 8028, 1144, -8165, -171, 8184, -807, -8089, 1773, 7876, -2718, -7551, 3623, 7114, -4480, -6576, 5271, 5940, -5989, -5217, 6618, 4416, -7154, -3550, 7583, 2628, -7904, -1668, 8106, 679, -8190, 319, 8149, -1317, -7989, 2294, 7707, -3240, -7310, 4138, 6800, -4976, -6188, 5738, 5479, -6416, -4687, 6994, 3820, -7469, -2895, 7827, 1921, -8067, -918, 8180, -103, -8169, 1122, 8027, -2127, -7762, 3099, 7372, -4025, -6868, 4887, 6252, -5676, -5537, 6373, 4732, -6972, -3851, 7458, 2905, -7828, -1913, 8069, 886, -8183, 154, 8163, -1196, -8011, 2218, 7726, -3208, -7317, 4144, 6784, -5016, -6141, 5805, 5393, -6500, -4556, 7087, 3640, -7558, -2664, 7902, 1639, -8115, -588, 8190, -478, -8129, 1535, 7928, -2569, -7594, 3560, 7128, -4493, -6541, 5349, 5839, -6116, -5037, 6776, 4144, -7323, -3181, 7741, 2158, -8027, -1099, 8171, 16, -8175, 1067, 8032, -2134, -7749, 3164, 7327, -4141, -6776, 5044, 6102, -5860, -5319, 6571, 4438, -7167, -3478, 7633, 2451, -7963, -1380, 8148, 281, -8187, 823, 8075, -1916, -7817, 2973, 7413, -3979, -6873, 4912, 6205, -5757, -5422, 6495, 4535, -7115, -3565, 7601, 2524, -7947, -1436, 8143, 318, -8188, 806, 8076, -1919, -7813, 2995, 7398, -4017, -6845, 4962, 6157, -5816, -5352, 6557, 4441, -7175, -3445, 7653, 2379, -7985, -1266, 8161, 126, -8179, 1017, 8036, -2143, -7737, 3227, 7283, -4251, -6686, 5191, 5954, -6031, -5105, 6750, 4151, -7337, -3114, 7777, 2012, -8063, -869, 8185, -295, -8145, 1452, 7937, -2584, -7569, 3663, 7045, -4671, -6378, 5582, 5578, -6383, -4664, 7051, 3650, -7577, -2561, 7944, 1416, -8149, -241, 8183, -942, -8048, 2105, 7742, -3228, -7275, 4282, 6652, -5250, -5890, 6106, 4999, -6836, -4004, 7419, 2919, -7846, -1773, 8105, 584, -8191, 616, 8100, -1807, -7835, 2958, 7399, -4049, -6803, 5052, 6056, -5948, -5178, 6712, 4183, -7333, -3097, 7792, 1939, -8081, -739, 8189, -482, -8119, 1691, 7865, -2866, -7438, 3977, 6842, -5003, -6093, 5915, 5205, -6698, -4199, 7328, 3096, -7795, -1922, 8084, 701, -8191, 535, 8109, -1763, -7843, 2951, 7395, -4074, -6777, 5102, 6000, -6016, -5085, 6790, 4049, -7409, -2919, 7854, 1717, -8117, -475, 8189, -781, -8070, 2019, 7759, -3213, -7266, 4330, 6598, -5348, -5774, 6238, 4809, -6983, -3730, 7559, 2558, -7957, -1325, 8161, 57, -8171, 1213, 7981, -2457, -7599, 3641, 7030, -4739, -6291, 5722, 5394, -6568, -4366, 7251, 3228, -7759, -2010, 8074, 739, -8191, 550, 8103, -1829, -7815, 3063, 7330, -4223, -6663, 5277, 5826, -6202, -4843, 6970, 3734, -7564, -2532, 7966, 1262, -8169, 40, 8161, -1345, -7947, 2615, 7528, -3821, -6916, 4929, 6124, -5914, -5175, 6744, 4089, -7404, -2897, 7870, 1627, -8133, -314, 8183, -1010, -8021, 2308, 7646, -3549, -7071, 4695, 6307, -5722, -5377, 6596, 4302, -7298, -3113, 7805, 1837, -8106, -513, 8189, -829, -8054, 2148, 7701, -3413, -7141, 4586, 6386, -5638, -5458)        
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L32C32_i
    );

    L32C33_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (2123, 8056, -820, -8190, -505, 8107, 1814, -7816, -3075, 7319, 4253, -6636, -5321, 5779, 6249, -4777, -7016, 3651, 7600, -2435, -7991, 1157, 8175, 148, -8152, -1449, 7920, 2710, -7490, -3902, 6869, 4992, -6077, -5957, 5132, 6769, -4061, -7413, 2888, 7868, -1647, -8129, 364, 8186, 924, -8041, -2190, 7696, 3398, -7164, -4522, 6454, 5532, -5589, -6408, 4586, 7123, -3475, -7666, 2279, 8021, -1031, -8182, -242, 8143, 1505, -7911, -2733, 7486, 3891, -6885, -4957, 6118, 5901, -5209, -6705, 4174, 7347, -3044, -7816, 1842, 8098, -600, -8191, -656, 8090, 1894, -7801, -3087, 7329, 4205, -6688, -5225, 5892, 6121, -4961, -6876, 3916, 7470, -2784, -7893, 1587, 8132, -358, -8187, -880, 8054, 2094, -7739, -3261, 7247, 4350, -6594, -5342, 5791, 6210, -4861, -6939, 3822, 7510, -2700, -7914, 1518, 8139, -305, -8186, -914, 8049, 2109, -7737, -3259, 7252, 4333, -6611, -5312, 5825, 6172, -4914, -6899, 3896, 7472, -2796, -7884, 1636, 8124, -444, -8190, -758, 8078, 1940, -7795, -3081, 7344, 4152, -6739, -5136, 5990, 6007, -5117, -6752, 4135, 7351, -3069, -7797, 1939, 8077, -772, -8190, -412, 8129, 1584, -7902, -2722, 7509, 3801, -6964, -4802, 6274, 5701, -5458, -6483, 4530, 7130, -3512, -7632, 2422, 7977, -1287, -8161, 125, 8178, 1035, -8032, -2175, 7723, 3267, -7261, -4295, 6654, 5233, -5916, -6068, 5061, 6780, -4108, -7358, 3074, 7789, -1983, -8067, 852, 8186, 291, -8146, -1429, 7946, 2536, -7593, -3594, 7093, 4578, -6458, -5475, 5698, 6264, -4832, -6933, 3873, 7467, -2843, -7860, 1759, 8101, -645, -8191, -481, 8124, 1595, -7907, -2678, 7539, 3708, -7033, -4670, 6395, 5541, -5641, -6310, 4782, 6959, -3838, -7480, 2823, 7862, -1760, -8101, 664, 8190, 441, -8131, -1537, 7923, 2602, -7574, -3621, 7088, 4570, -6476, -5439, 5747, 6206, -4919, -6864, 4003, 7396, -3019, -7799, 1981, 8061, -912, -8183, -174, 8159, 1252, -7995, -2310, 7689, 3323, -7252, -4279, 6688, 5157, -6011, -5947, 5230, 6632, -4363, -7204, 3420, 7650, -2422, -7967, 1383, 8146, -324, -8189, -741, 8092, 1789, -7861, -2808, 7497, 3776, -7010, -4682, 6405, 5506, -5697, -6240, 4894, 6868, -4014, -7383, 3067, 7775, -2073, -8041, 1046, 8174, -5, -8175, -1037, 8042, 2058, -7782, -3046, 7395, 3982, -6892, -4854, 6278, 5645, -5567, -6348, 4767, 6947, -3895, -7437, 2961, 7807, -1984, -8056, 975, 8177, 45, -8173, -1064, 8039, 2064, -7784, -3032, 7406, 3949, -6918, -4807, 6323, 5587, -5634, -6283, 4858, 6880, -4012, -7375, 3105, 7755, -2155, -8020, 1173, 8163, -176, -8185, -824, 8084, 1807, -7865, -2765, 7528, 3677, -7083, -4537, 6533, 5326, -5890, -6038, 5161, 6659, -4360, -7185, 3495, 7604, -2584, -7914, 1635, 8109, -666, -8190, -313, 8151, 1283, -8000, -2236, 7733, 3153, -7360, -4026, 6882, 4840, -6311, -5586, 5651, 6251, -4916, -6831, 4111, 7313, -3254, -7695, 2352, 7970, -1420, -8137, 470, 8190, 484, -8135, -1431, 7968, 2355, -7696, -3248, 7319, 4094, -6846, -4885, 6282, 5609, -5637, -6258, 4917, 6822, -4135, -7297, 3298, 7673, -2422, -7951, 1514, 8122, -590, -8191, -342, 8151, 1266, -8008, -2174, 7761, 3051, -7418, -3889, 6978, 4674, -6453, -5400, 5846, 6055, -5168, -6635, 4425, 7129, -3629, -7535, 2789, 7844, -1917, -8058, 1021, 8171, -116, -8185, -790, 8096, 1683, -7912, -2556, 7629, 3394, -7257, -4192, 6796, 4936, -6257, -5621, 5642, 6236, -4963, -6778, 4224, 7236, -3439, -7610, 2613, 7892, -1760, -8084, 886, 8178, -6, -8180, -875, 8085, 1742, -7899, -2590, 7621, 3404, -7258, -4179, 6812, 4904, -6291, -5574, 5698, 6177, -5044, -6712, 4333, 7169, -3577, -7548, 2781, 7839, -1958, -8046, 1112, 8162, -259, -8190, -598, 8126, 1445, -7977, -2276, 7739, 3079, -7420, -3850, 7021, 4575, -6549, -5252, 6006, 5870, -5403, -6427, 4742, 6912, -4034, -7327, 3284, 7661, -2502, -7917, 1695, 8089, -873, -8179, 43, 8182, 785, -8104, -1605, 7941, 2404, -7700, -3180, 7379, 3920, -6987, -4621, 6523, 5272, -5998, -5872, 5412, 6409, -4775, -6885, 4091, 7290, -3370, -7624, 2615, 7881, -1839, -8063, 1045, 8165, -244, -8190, -559, 8134, 1354, -8003, -2136, 7794, 2893, -7514, -3624, 7161, 4317, -6744, -4971, 6263, 5574, -5726, -6126, 5136, 6619, -4502, -7052, 3826, 7417, -3118, -7715, 2381, 7941, -1627, -8097, 857, 8177, -84, -8186, -691, 8120, 1456, -7984, -2208, 7775, 2937, -7501, -3640, 7159, 4308, -6758, -4939, 6297, 5524, -5785, -6062, 5222, 6545, -4617, -6972, 3973, 7338, -3298, -7642, 2595, 7879, -1874, -8052, 1137, 8155, -394, -8191, -353, 8158, 1093, -8060, -1824, 7894, 2537, -7666, -3229, 7374, 3892, -7026, -4523, 6619, 5115, -6163, -5667, 5656, 6170, -5108, -6625, 4518, 7025, -3897, -7371, 3245, 7656, -2570, -7883, 1876, 8047, -1171, -8151, 456, 8190, 258, -8168, -971, 8083, 1672, -7939, -2362, 7733, 3029, -7473, -3675, 7155, 4290, -6787, -4874, 6368, 5418, -5906, -5924, 5399, 6383, -4857, -6797, 4279, 7159, -3673, -7471, 3041, 7726, -2391, -7929, 1724, 8072, -1048, -8161, 364, 8190, 318, -8165, -999, 8081, 1669, -7944, -2327, 7750, 2967, -7506, -3586, 7210, 4177, -6869, -4741, 6480, 5270, -6050, -5764, 5580, 6217, -5076, -6630, 4538, 6996, -3974, -7318, 3383, 7589, -2774, -7813, 2147, 7984, -1509, -8105, 862, 8173, -213, -8191, -438, 8155, 1082, -8071, -1720, 7934, 2343, -7751, -2952, 7519, 3540, -7243, -4106, 6922, 4644, -6562, -5155, 6161, 5631, -5727, -6074, 5258, 6478, -4760, -6844, 4235, 7168, -3687, -7450, 3118, 7687, -2535, -7880, 1936, 8026, -1330, -8127, 716, 8180, -102, -8189, -513, 8150, 1122, -8067, -1724, 7937, 2314, -7767, -2891, 7552, 3448, -7298, -3987, 7003, 4501, -6674, -4991, 6308, 5451, -5911, -5883, 5481, 6281, -5027, -6646, 4545, 6973, -4043, -7266, 3519, 7517, -2981, -7732, 2427, 7904, -1864, -8038, 1292, 8129, -716, -8180, 137, 8189, 439, -8159, -1013, 8087, 1578, -7978, -2137, 7828, 2681, -7643, -3212, 7419, 3724, -7163, -4220, 6871, 4691, -6550, -5141, 6197, 5564, -5818, -5961, 5412, 6328, -4983, -6666, 4532, 6971, -4063, -7246, 3575, 7485, -3074, -7691, 2560, 7861, -2038, -7997, 1506, 8096, -972, -8161, 433, 8189, 105, -8183, -642, 8140, 1172, -8065, -1698, 7953, 2213, -7811, -2719, 7634, 3210, -7429, -3688, 7191, 4148, -6927, -4591, 6634, 5012, -6316, -5413, 5973, 5790, -5609, -6144, 5221, 6471, -4817, -6773, 4393, 7046, -3955, -7293, 3502, 7509, -3039, -7697, 2564, 7854, -2083, -7983, 1593, 8079, -1102, -8147, 606, 8183, -111, -8190, -384, 8166, 874, -8115, -1361, 8032, 1840, -7924, -2312, 7785, 2773, -7622, -3224, 7431, 3661, -7217, -4085, 6977, 4492, -6716, -4884, 6431, 5256, -6128, -5611, 5803, 5944, -5462, -6259, 5103, 6550, -4730, -6820, 4341, 7065, -3942, -7289, 3530, 7487, -3110, -7663, 2680, 7811, -2245, -7937, 1802, 8037, -1358, -8113, 910, 8162, -462, -8188, 13, 8188, 433, -8165, -877, 8117, 1316, -8047, -1750, 7952, 2176, -7836, -2596, 7696, 3005, -7538, -3406, 7356, 3794, -7157, -4172, 6937, 4534, -6701, -4885, 6445, 5220, -6175, -5540, 5888, 5843, -5588, -6131, 5273, 6400, -4947, -6653, 4608, 6886, -4260, -7102, 3901, 7297, -3536, -7476, 3161, 7632, -2782, -7771, 2396, 7889, -2007, -7989, 1613, 8067, -1219, -8128, 822, 8167, -427, -8188, 31, 8189, 362, -8172, -755, 8135, 1142, -8082, -1526, 8009, 1904, -7920, -2277, 7812, 2642, -7690, -3002, 7549, 3351, -7395, -3694, 7224, 4025, -7040, -4348, 6840, 4659, -6629, -4961, 6404, 5249, -6169, -5527, 5920, 5791, -5662, -6044, 5393, 6282, -5116, -6509, 4829, 6719, -4536, -6919, 4234, 7102, -3927, -7272, 3612, 7427, -3294, -7569, 2970, 7694, -2644, -7808, 2312, 7904, -1981, -7988, 1645, 8056, -1310, -8112, 973, 8151, -638, -8178, 301, 8189, 32, -8189, -365, 8173, 695, -8146, -1023, 8104, 1346, -8052, -1667, 7985, 1982, -7907, -2294, 7816, 2599, -7716, -2900, 7602, 3194, -7480, -3483, 7345, 3763, -7203, -4038, 7048, 4304, -6887, -4564, 6714, 4815, -6536, -5059, 6347, 5293, -6152, -5521, 5949, 5737, -5740, -5947, 5524, 6146, -5303, -6338, 5075, 6518, -4843, -6692, 4605, 6853, -4365, -7008, 4118, 7150, -3870, -7286, 3617, 7409, -3363, -7526, 3105, 7631, -2847, -7728, 2585, 7814, -2324, -7893, 2060, 7960, -1797, -8020, 1533, 8070, -1270, -8112, 1005, 8144, -743, -8169, 480, 8183, -221, -8191, -39, 8189, 296, -8181, -552, 8162, 804, -8138, -1056, 8105, 1303, -8066, -1549, 8018, 1790, -7966, -2029, 7904, 2264, -7838, -2496, 7764, 2723, -7685, -2947, 7599, 3166, -7508, -3382, 7411, 3592, -7310, -3800, 7202, 4001, -7091, -4200, 6974, 4391, -6854, -4580, 6728, 4762, -6599, -4941, 6466, 5114, -6330, -5283, 6189, 5445, -6047, -5604, 5900, 5756, -5753, -5905, 5600, 6047, -5448, -6186, 5291, 6318, -5134, -6447, 4973, 6568, -4813, -6687, 4649, 6799, -4485, -6908, 4319, 7010, -4154, -7109, 3986, 7201, -3819, -7291, 3649, 7374, -3482, -7454, 3312, 7528, -3143, -7599, 2973, 7664, -2805, -7726, 2636, 7783, -2469, -7837, 2300, 7885, -2134, -7931, 1966, 7971, -1802, -8009, 1636, 8042, -1473, -8072, 1310, 8098, -1149, -8121, 988, 8140, -830, -8157, 672, 8169, -517, -8180, 362, 8186, -210, -8190, 58, 8190, 91, -8190, -239, 8185, 384, -8179, -529, 8169, 670, -8158, -811, 8143, 949, -8128, -1086, 8109, 1219, -8090, -1352, 8067, 1481, -8044, -1610, 8018, 1735, -7992, -1860, 7962, 1981, -7933, -2102, 7901, 2218, -7869, -2334, 7834, 2446, -7800, -2558, 7763, 2666, -7727, -2774, 7688, 2878, -7650, -2981, 7609, 3080, -7570, -3179, 7528, 3274, -7488, -3369, 7445, 3460, -7403, -3551, 7360, 3637, -7318, -3724, 7274, 3807, -7231, -3889, 7187, 3968, -7144, -4046, 7100, 4121, -7057, -4195, 7013, 4266, -6971, -4337, 6927, 4404, -6885, -4471, 6842, 4534, -6801, -4597, 6758, 4657, -6718, -4717, 6676, 4773, -6637, -4829, 6596, 4881, -6558, -4934, 6519, 4983, -6482, -5033, 6444, 5079, -6409, -5125, 6372, 5167, -6338, -5210, 6303, 5250, -6271, -5290, 6238, 5326, -6207, -5363, 6176, 5397, -6147, -5431, 6118, 5461, -6091, -5492, 6064, 5520, -6039, -5548, 6014, 5573, -5991, -5599, 5968, 5621, -5947, -5644, 5926, 5663, -5908, -5684, 5889, 5701, -5874, -5718, 5857, 5733, -5844, -5748, 5829, 5760, -5818, -5772, 5806, 5781, -5798, -5792, 5788, 5798, -5782, -5806, 5775, 5810, -5771, -5816, 5767, 5818, -5765, -5820, 5763, 5820, -5764, -5820, 5764, 5817, -5768, -5815, 5771, 5810, -5777, -5805, 5782, 5797, -5790, -5790, 5798, 5780, -5809, -5771, 5819, 5758, -5832, -5746, 5845, 5730, -5860, -5716, 5875, 5698, -5893, -5681, 5910, 5661, -5930, -5641, 5949, 5618, -5972, -5595, 5993, 5570, -6018, -5544, 6042, 5516, -6068, -5488, 6094, 5457, -6123, -5426, 6151, 5392, -6181, -5358, 6211, 5321, -6243, -5284, 6275, 5244, -6309, -5204, 6342, 5161, -6378, -5118, 6413, 5072, -6450, -5026, 6486, 4976, -6525, -4927, 6563, 4874, -6603, -4821, 6642, 4764, -6683, -4708, 6723, 4648, -6765, -4588, 6806, 4525, -6849, -4461, 6890, 4394, -6934, -4327, 6976, 4256, -7020, -4185, 7063, 4110, -7107, -4035, 7150, 3956, -7194, -3878, 7237, 3795, -7281, -3712, 7323, 3625, -7367, -3538, 7408, 3447, -7452, -3356, 7493, 3261, -7535, -3165, 7575, 3066, -7616, -2966, 7654, 2863, -7694, -2759, 7731, 2651, -7769, -2543, 7804, 2430, -7840, -2318, 7873, 2201, -7906, -2084, 7936, 1964, -7967, -1843, 7995, 1717, -8023, -1592, 8047, 1463, -8071, -1333, 8092, 1200, -8113, -1066, 8129, 929, -8146, -791, 8159, 650, -8171, -508, 8179, 363, -8186, -218, 8189, 69, -8191, 80, 8189, -232, -8186, 384, 8177, -540, -8168, 695, 8154, -853, -8138, 1011, 8117, -1173, -8095, 1333, 8067, -1497, -8038, 1660, 8003, -1826, -7966, 1990, 7924, -2158, -7879, 2324, 7828, -2493, -7776, 2660, 7717, -2830, -7656, 2998, 7588, -3168, -7518, 3336, 7442, -3506, -7363, 3674, 7277, -3843, -7189, 4010, 7094, -4178, -6996, 4343, 6892, -4509, -6784, 4672, 6670, -4836, -6552, 4996, 6428, -5157, -6300, 5313, 6166, -5470, -6028, 5622, 5883, -5774, -5736, 5922, 5581, -6068, -5423, 6210, 5258, -6350, -5090, 6485, 4915, -6618, -4737, 6746, 4552, -6871, -4365, 6991, 4170, -7107, -3973, 7218, 3769, -7325, -3563, 7425, 3351, -7522, -3136, 7611, 2914, -7697, -2691, 7775, 2462, -7848, -2231, 7913, 1994, -7974, -1756, 8026, 1513, -8073, -1268, 8110, 1019, -8143, -769, 8165, 515, -8182, -260, 8189, 1, -8191, 257, 8181, -519, -8166, 780, 8140, -1044, -8107, 1307, 8063, -1572, -8012, 1835, 7951, -2099, -7882, 2361, 7802, -2624, -7715, 2884, 7616, -3144, -7510, 3399, 7392, -3655, -7267, 3905, 7130, -4155, -6986, 4399, 6830, -4641, -6667, 4876, 6493, -5109, -6311, 5334, 6118, -5556, -5918, 5770, 5707, -5979, -5489, 6180, 5260, -6375, -5025, 6561, 4779, -6741, -4527, 6910, 4266, -7072, -3999, 7223, 3723, -7366, -3441, 7498, 3152, -7620, -2857, 7730, 2555, -7831, -2250, 7918, 1937, -7996, -1621, 8059, 1299, -8112, -976, 8150, 647, -8177, -317, 8189, -16, -8189, 350, 8174, -687, -8147, 1022, 8104, -1359, -8048, 1694, 7976, -2029, -7892, 2360, 7791, -2691, -7678, 3017, 7548, -3340, -7406, 3658, 7248, -3971, -7077, 4277, 6890, -4579, -6691, 4871, 6476, -5157, -6249, 5432, 6007, -5700, -5754, 5956, 5487, -6203, -5209, 6437, 4917, -6661, -4616, 6870, 4301, -7067, -3979, 7249, 3644, -7418, -3302, 7570, 2950, -7708, -2591, 7829, 2223, -7934, -1850, 8020, 1470, -8091, -1087, 8142, 697, -8176, -307, 8190, -89, -8187, 483, 8162, -881, -8120, 1276, 8057, -1671, -7976, 2063, 7873, -2452, -7753, 2836, 7611, -3216, -7451, 3588, 7270, -3954, -7072, 4310, 6853, -4658, -6618, 4994, 6362, -5320, -6091, 5631, 5800, -5931, -5495, 6214, 5172, -6484, -4836, 6735, 4483, -6971, -4118, 7186, 3739, -7384, -3349, 7561, 2947, -7719, -2536, 7853, 2115, -7968, -1688, 8057, 1252, -8126, -813, 8169, 368, -8190, 78, 8185, -527, -8157, 974, 8102, -1423, -8025, 1866, 7920, -2308, -7792, 2742, 7638, -3171, -7461, 3590, 7258, -4001, -7032, 4398, 6781, -4785, -6510, 5156, 6214, -5513, -5898, 5851, 5560, -6173, -5204, 6473, 4827, -6755, -4435, 7013, 4024, -7250, -3599, 7460, 3159, -7648, -2708, 7807, 2244, -7941, -1772, 8046, 1290, -8124, -804, 8171, 312, -8191, 182, 8179, -678, -8139, 1172, 8067, -1665, -7966, 2152, 7833, -2634, -7672, 3106, 7479, -3569, -7259, 4019, 7008, -4456, -6731, 4876, 6425, -5279, -6095, 5662, 5737, -6025, -5357, 6363, 4952, -6679, -4528, 6966, 4083, -7228, -3621, 7460, 3140, -7663, -2647, 7833, 2139, -7972, -1623, 8077, 1096, -8149, -564, 8185, 27, -8188, 510, 8153, -1049, -8085, 1583, 7979, -2114, -7840, 2635, 7663, -3148, -7453, 3646, 7207, -4132, -6930, 4598, 6619, -5047, -6278, 5472, 5905, -5875, -5505, 6249, 5077, -6598, -4625, 6915, 4148, -7202, -3652, 7453, 3135, -7672, -2604, 7852, 2056, -7996, -1498, 8100, 930, -8166, -357, 8190, -222, -8176, 799, 8118, -1376, -8021, 1945, 7882, -2508, -7704, 3058, 7483, -3597, -7226, 4116, 6928, -4617, -6595, 5093, 6225, -5546, -5823, 5969, 5387, -6363, -4922, 6723, 4428, -7049, -3911, 7336, 3369, -7586, -2808, 7793, 2229, -7960, -1638, 8081, 1034, -8159, -425, 8190, -191, -8176, 805, 8115, -1418, -8009, 2023, 7854, -2620, -7656, 3201, 7411, -3768, -7124, 4312, 6793, -4834, -6423, 5327, 6011, -5792, -5565, 6221, 5082, -6616, -4569, 6971, 4025, -7286, -3457, 7555, 2865, -7781, -2255, 7957, 1627, -8086, -990, 8163, 343, -8191, 306, 8166, -957, -8091, 1601, 7962, -2239, -7784, 2862, 7553, -3470, -7274, 4056, 6946, -4618, -6573, 5150, 6154, -5651, -5696, 6114, 5196, -6539, -4662, 6920, 4094, -7257, -3498, 7544, 2875, -7782, -2233, 7966, 1573, -8097, -901, 8171, 220, -8191, 463, 8151, -1146, -8056, 1821, 7902, -2486, -7694, 3134, 7428, -3763, -7111, 4364, 6739, -4938, -6320, 5475, 5853, -5975, -5343, 6431, 4791, -6843, -4204, 7204, 3583, -7514, -2935, 7766, 2262, -7963, -1573, 8099, 867, -8175, -156, 8188, -561, -8140, 1272, 8027, -1978, -7855, 2668, 7618, -3341, -7324, 3988, 6970, -4607, -6562, 5189, 6100, -5733, -5590, 6231, 5032, -6682, -4434, 7079, 3798, -7421, -3131, 7702, 2435, -7923, -1720, 8078, 986, -8168, -245, 8190, -501, -8145, 1244, 8030, -1979, -7850, 2698, 7601, -3398, -7290, 4068, 6913, -4707, -6479, 5306, 5987, -5862, -5443, 6367, 4850, -6820, -4215, 7212, 3540, -7545, -2834, 7809, 2099, -8008, -1347, 8134, 579, -8189, 195, 8170, -970, -8079, 1736, 7913, -2490, -7677, 3221, 7368, -3926, -6993, 4595, 6551, -5225, -6050, 5806, 5490, -6337, -4879, 6807, 4220, -7217, -3521, 7558, 2785, -7830, -2024, 8026, 1240, -8148, -444, 8190, -360, -8156, 1160, 8041, -1953, -7850, 2726, 7579, -3476, -7236, 4192, 6820, -4870, -6337, 5499, 5788, -6078, -5182, 6594, 4522, -7048, -3816, 7430, 3069, -7739, -2291, 7969, 1486, -8120, -667, 8187, -164, -8171, 992, 8069, -1814, -7886, 2616, 7618, -3395, -7272, 4138, 6847, -4841, -6351, 5493, 5785, -6090, -5158, 6621, 4473, -7084, -3741, 7471, 2965, -7779, -2158, 8003, 1323, -8142, -475, 8190, -382, -8151, 1235, 8021, -2078, -7803, 2898, 7497, -3689, -7109, 4439, 6639, -5142, -6095, 5787, 5480, -6371, -4804, 6881, 4069, -7316, -3289, 7666, 2468, -7932, -1619, 8104, 748, -8186, 132, 8170, -1014, -8062, 1884, 7857, -2735, -7562, 3554, 7175, -4335, -6704, 5064, 6152, -5736, -5526, 6339, 4832, -6869, -4080, 7316, 3276, -7677, -2432, 7943, 1555, -8116, -660, 8188, -247, -8162, 1151, 8033, -2044, -7806, 2912, 7481, -3747, -7064, 4535, 6556, -5270, -5966, 5938, 5299, -6534, -4565, 7047, 3770, -7473, -2927, 7803, 2044, -8035, -1135, 8163, 207, -8187, 723, 8104, -1647, -7917, 2550, 7625, -3423, -7234, 4250, 6746, -5026, -6169, 5734, 5508, -6370, -4775, 6920, 3975, -7380, -3122, 7741, 2223, -8000, -1295, 8149, 346, -8190, 607, 8119, -1556, -7938, 2484, 7646, -3381, -7250, 4231, 6752, -5026, -6161, 5751, 5482, -6399, -4727, 6957, 3903, -7420, -3024, 7778, 2099, -8029, -1145, 8164, 170, -8185, 806, 8088, -1774, -7877, 2717, 7550, -3624, -7115, 4479, 6575, -5272, -5941, 5988, 5216, -6619, -4417, 7153, 3549, -7584, -2629, 7903, 1667, -8107, -680, 8189, -320, -8150, 1316, 7988, -2295, -7708, 3239, 7309, -4139, -6801, 4975, 6187, -5739, -5480, 6415, 4686, -6995, -3821, 7468, 2894, -7828, -1922, 8066, 917, -8181, 102, 8168, -1123, -8028, 2126, 7761, -3100, -7373, 4024, 6867, -4888, -6253, 5675, 5536, -6374, -4733, 6971, 3850, -7459, -2906, 7827, 1912, -8070, -887, 8182, -155, -8164, 1195, 8010, -2219, -7727, 3207, 7316, -4145, -6785, 5015, 6140, -5806, -5394, 6499, 4555, -7088, -3641, 7557, 2663, -7903, -1640, 8114, 587, -8191, 477, 8128, -1536, -7929, 2568, 7593, -3561, -7129, 4492, 6540, -5350, -5840, 6115, 5036, -6777, -4145, 7322, 3180, -7742, -2159, 8026, 1098, -8172, -17, 8174, -1068, -8033, 2133, 7748, -3165, -7328, 4140, 6775, -5045, -6103, 5859, 5318, -6572, -4439, 7166, 3477, -7634, -2452, 7962, 1379, -8149, -282, 8186, -824, -8076, 1915, 7816, -2974, -7414, 3978, 6872, -4913, -6206, 5756, 5421, -6496, -4536, 7114, 3564, -7602, -2525, 7946, 1435, -8144, -319, 8187, -807, -8077, 1918, 7812, -2996, -7399, 4016, 6844, -4963, -6158, 5815, 5351, -6558, -4442, 7174, 3444, -7654, -2380, 7984, 1265, -8162, -127, 8178, -1018, -8037, 2142, 7736, -3228, -7284, 4250, 6685, -5192, -5955, 6030, 5104, -6751, -4152, 7336, 3113, -7778, -2013, 8062, 868, -8186, 294, 8144, -1453, -7938, 2583, 7568, -3664, -7046, 4670, 6377, -5583, -5579, 6382, 4663, -7052, -3651, 7576, 2560, -7945, -1417, 8148, 240, -8184, 941, 8047, -2106, -7743, 3227, 7274, -4283, -6653, 5249, 5889, -6107, -5000, 6835, 4003, -7420, -2920, 7845, 1772, -8106, -585, 8190, -617, -8101, 1806, 7834, -2959, -7400, 4048, 6802, -5053, -6057, 5947, 5177, -6713, -4184, 7332, 3096, -7793, -1940, 8080, 738, -8190, 481, 8118, -1692, -7866, 2865, 7437, -3978, -6843, 5002, 6092, -5916, -5206, 6697, 4198, -7329, -3097, 7794, 1921, -8085, -702, 8190, -536, -8110, 1762, 7842, -2952, -7396, 4073, 6776, -5103, -6001, 6015, 5084, -6791, -4050, 7408, 2918, -7855, -1718, 8116, 474, -8190, 780, 8069, -2020, -7760, 3212, 7265, -4331, -6599, 5347, 5773, -6239, -4810, 6982, 3729, -7560, -2559, 7956, 1324, -8162, -58, 8170, -1214, -7982, 2456, 7598, -3642, -7031, 4738, 6290, -5723, -5395, 6567, 4365, -7252, -3229, 7758, 2009, -8075, -740, 8190, -551, -8104, 1828, 7814, -3064, -7331, 4222, 6662, -5278, -5827, 6201, 4842, -6971, -3735, 7563, 2531, -7967, -1263, 8168, -41, -8162, 1344, 7946, -2616, -7529, 3820, 6915, -4930, -6125, 5913, 5174, -6745, -4090, 7403, 2896, -7871, -1628, 8132, 313, -8184, 1009, 8020, -2309, -7647, 3548, 7070, -4696, -6308, 5721, 5376, -6597, -4303, 7297, 3112, -7806, -1838, 8105, 512, -8190, 828, 8053, -2149, -7702, 3412, 7140, -4587, -6387, 5637, 5457)         
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L32C33_i
    );

process(Clk_96, Ce_F6 , TI , LG  )
    variable count: integer := 0;
    variable guard: boolean := False;
begin
    if TI = '1' then    
        adress <= "11";
    elsif rising_edge(clk_96) then         
            if LG = '0' and guard = False  then                          
                 guard := True;
                 adress <= adress +1;                                    
                if adress = "11" then
                   adress <= "00";
                end if;
            elsif LG = '1' then 
               guard := False;
            end if;     
    end if;                                      
end process;

    pft_adress <= PFT & adress ;
process(PFT_adress, Rom_cos_L15_i, Rom_cos_L15�31_i, Rom_cos_L15�32_i, Rom_cos_L15�33_i, Rom_cos_L21_i, Rom_cos_L21C31_i, Rom_cos_L21C32_i, Rom_cos_L21C33_i, Rom_cos_L32_i, Rom_cos_L32C31_i, Rom_cos_L32C32_i, Rom_cos_L32C33_i)
begin
  if  pft_adress = "0110000000" or pft_adress = "0110001100" then
        Rom_cos_i <= Rom_cos_L15_i;
    elsif pft_adress = "0110000100" or pft_adress = "0110001000" or pft_adress = "0110011000" or pft_adress = "0110011100" or pft_adress = "0111000100" or pft_adress = "0111001000" or pft_adress = "0111011000" or pft_adress = "0111011100" then
        Rom_cos_i <= Rom_cos_L15�31_i;
    elsif pft_adress = "0110000101" or pft_adress = "0110001001" or pft_adress = "0110011001" or pft_adress = "0110011101" or pft_adress = "0111000101" or pft_adress = "0111001001" or pft_adress = "0111011001" or pft_adress = "0111011101" then
        Rom_cos_i <= Rom_cos_L15�32_i;
    elsif pft_adress = "0110000110" or pft_adress = "0110001010" or pft_adress = "0110011010" or pft_adress = "0110011110" or pft_adress = "0111000110" or pft_adress = "0111001010" or pft_adress = "0111011010" or pft_adress = "0111011110" then
        Rom_cos_i <= Rom_cos_L15�33_i;
    elsif pft_adress = "0100000000" or pft_adress = "0100001100" then
        Rom_cos_i <= Rom_cos_L21_i;
    elsif pft_adress = "0100000100" or pft_adress = "0100001000" or pft_adress = "0100011000" or pft_adress = "0100011100" or pft_adress = "0101000100" or pft_adress = "0101001000" or pft_adress = "0101011000" or pft_adress = "0101011100" then
        Rom_cos_i <= Rom_cos_L21C31_i;
    elsif pft_adress = "0100000101" or pft_adress = "0100001001" or pft_adress = "0100011001" or pft_adress = "0100011101" or pft_adress = "0101000101" or pft_adress = "0101001001" or pft_adress = "0101011001" or pft_adress = "0101011101" then
        Rom_cos_i <= Rom_cos_L21C32_i;
    elsif pft_adress = "0100000110" or pft_adress = "0100001010" or pft_adress = "0100011010" or pft_adress = "0100011110" or pft_adress = "0101000110" or pft_adress = "0101001010" or pft_adress = "0101011010" or pft_adress = "0101011110" then
        Rom_cos_i <= Rom_cos_L21C33_i;
    elsif pft_adress = "0010000000" or pft_adress = "0010001100" then
        Rom_cos_i <= Rom_cos_L32_i;
    elsif pft_adress = "0010000100" or pft_adress = "0010001000" or pft_adress = "0010011000" or pft_adress = "0010011100" or pft_adress = "0011000100" or pft_adress = "0011001000" or pft_adress = "0011011000" or pft_adress = "0011011100" then
        Rom_cos_i <= Rom_cos_L32C31_i;
    elsif pft_adress = "0010000101" or pft_adress = "0010001001" or pft_adress = "0010011001" or pft_adress = "0010011101" or pft_adress = "0011000101" or pft_adress = "0011001001" or pft_adress = "0011011001" or pft_adress = "0011011101" then
        Rom_cos_i <= Rom_cos_L32C32_i;
    elsif pft_adress = "0010000110" or pft_adress = "0010001010" or pft_adress = "0010011010" or pft_adress = "0010011110" or pft_adress = "0011000110" or pft_adress = "0011001010" or pft_adress = "0011011010" or pft_adress = "0011011110" then
        Rom_cos_i <= Rom_cos_L32C33_i;
    end if; 
 end process;

process (Clk_96, Ce_F6, EN, Rom_cos_i )
begin
         
    if EN = '1' then
       Rom_cos <= conv_std_logic_vector(Rom_cos_i- magic, data_rom);
    else
       Rom_cos <=(others => '0');
    end if;     
end process;end Behavioral;
