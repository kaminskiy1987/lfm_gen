
--������������� �� ������------ �� �������--------
library IEEE;
	use IEEE.STD_LOGIC_1164.ALL;
	Use ieee.std_logic_arith.all;
	Use ieee.std_logic_unsigned.all;
	USE ieee.math_real.all;
	USE std.textio.ALL;
	USE IEEE.std_logic_textio.ALL;

library elementary;
	use elementary.s274types_pkg.all;
	use elementary.utility.all;
	use elementary.all;
    
entity MUX_signal_type4 is
       generic (
	
	   data_pft: integer := 6;
		data_ppz : integer := 5;
		pft_widht : integer:= 6;
		pft_code : int_array := (10,27);
		data_rom : integer := 12
				);
	Port(
		Clk_96 : in std_logic;
		Ce_F6 : in std_logic;
		En : in std_logic;      
		OD : in std_logic;		
	        LG : in std_logic;		
	        TI : in std_logic;
		PFT : in std_logic_vector (7 downto 0);		
		Sign_LCHM : in std_logic;
		Rom_cos : out std_logic_vector (13 downto 0)		
	);

end MUX_signal_type4;

architecture Behavioral of MUX_signal_type4 is

	signal P2_PFT : std_logic_vector(7 downto 0) := (others => '0');
    signal PFT_adress : std_logic_vector(9 downto 0) := (others => '0');
	signal Rom_cos_i : integer;
	signal adress : std_logic_vector(1 downto 0);  
	signal Rom_cos_L15_i : integer;
	signal Rom_cos_L15�31_i : integer;
	signal Rom_cos_L15�32_i : integer;
	signal Rom_cos_L15�33_i : integer;
	signal Rom_cos_L21_i : integer;
	signal Rom_cos_L21C31_i : integer;
	signal Rom_cos_L21C32_i : integer;
	signal Rom_cos_L21C33_i : integer;
	signal Rom_cos_L32_i : integer;
	signal Rom_cos_L32C31_i : integer;
	signal Rom_cos_L32C32_i : integer;
	signal Rom_cos_L32C33_i : integer;
	signal Rom_cos_L40_i : integer;
	signal Rom_cos_L40C31_i : integer;
	signal Rom_cos_L40C32_i : integer;
	signal Rom_cos_L40C33_i : integer;
begin

    L15_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-5300, 4212, 8004, 919, -7418, -5663, 3801, 8088, 1349, -7232, -5943, 3463, 8137, 1683, -7075, -6148, 3202, 8163, 1925, -6957, -6285, 3025, 8175, 2075, -6884, -6360, 2933, 8180, 2135, -6861, -6375, 2927, 8179, 2105, -6888, -6332, 3008, 8173, 1984, -6964, -6228, 3175, 8158, 1773, -7085, -6060, 3425, 8126, 1469, -7245, -5821, 3754, 8069, 1070, -7432, -5503, 4156, 7974, 577, -7634, -5096, 4622, 7824, -12, -7833, -4591, 5139, 7602, -694, -8009, -3978, 5693, 7289, -1462, -8138, -3250, 6260, 6862, -2306, -8191, -2400, 6815, 6304, -3211, -8139, -1430, 7325, 5594, -4152, -7948, -346, 7753, 4719, -5097, -7586, 837, 8056, 3672, -6006, -7024, 2093, 8188, 2454, -6829, -6236, 3382, 8103, 1081, -7510, -5207, 4654, 7756, -416, -7984, -3935, 5844, 7109, -1990, -8188, -2437, 6874, 6140, -3573, -8060, -749, 7659, 4841, -5078, -7547, 1064, 8113, 3235, -6402, -6618, 2912, 8152, 1372, -7433, -5267, 4679, 7710, -661, -8056, -3525, 6228, 6749, -2741, -8165, -1465, 7412, 5270, -4713, -7682, 789, 8085, 3325, -6397, -6571, 3070, 8122, 1028, -7607, -4853, 5171, 7444, -1449, -8169, -2623, 6864, 6032, -3875, -7951, -54, 7925, 3954, -5984, -6890, 2610, 8166, 1373, -7499, -5019, 5064, 7471, -1453, -8174, -2485, 6980, 5834, -4186, -7837, 445, 8050, 3381, -6446, -6436, 3403, 8042, 385, -7863, -4076, 5954, 6860, -2754, -8144, -1033, 7665, 4582, -5548, -7143, 2258, 8181, 1494, -7499, -4921, 5254, 7313, -1933, -8191, -1774, 7390, 5104, -5095, -7394, 1782, 8190, 1873, -7358, -5145, 5075, 7392, -1810, -8191, -1796, 7402, 5041, -5199, -7312, 2013, 8187, 1539, -7522, -4791, 5456, 7139, -2391, -8165, -1102, 7695, 4379, -5835, -6855, 2933, 8094, 477, -7895, -3792, 6307, 6427, -3627, -7938, 330, 8075, 3008, -6835, -5824, 4443, 7645, -1317, -8184, -2017, 7364, 5003, -5341, -7160, 2456, 8147, 810, -7825, -3935, 6257, 6422, -3711, -7892, 595, 8126, 2598, -7109, -5381, 5008, 7331, -2160, -8170, -1001, 7784, 3997, -6250, -6393, 3805, 7845, -821, -8158, -2270, 7300, 5021, -5413, -7054, 2772, 8089, 240, -8001, -3207, 6815, 5721, -4710, -7452, 1980, 8175, 999, -7814, -3834, 6426, 6153, -4212, -7667, 1465, 8190, 1453, -7675, -4177, 6197, 6363, -3959, -7754, 1243, 8188, 1609, -7631, -4255, 6159, 6378, -3967, -7741, 1318, 8190, 1469, -7693, -4074, 6317, 6201, -4235, -7621, 1689, 8184, 1030, -7844, -3623, 6649, 5808, -4747, -7361, 2346, 8124, 287, -8033, -2878, 7107, 5156, -5460, -6898, 3266, 7933, -759, -8174, -1812, 7606, 4188, -6302, -6148, 4396, 7506, -2085, -8148, -411, 8022, 2853, -7157, -5021, 5641, 6718, -3627, -7804, 1300, 8190, 1127, -7858, -3443, 6847, 5448, -5258, -6979, 3233, 7913, -952, -8188, -1395, 7790, 3612, -6766, -5528, 5206, 6991, -3249, -7899, 1048, 8190, 1216, -7856, -3376, 6931, 5268, -5498, -6761, 3670, 7749, -1591, -8176, -591, 8019, 2715, -7303, -4637, 6087, 6227, -4466, -7388, 2555, 8046, -490, -8172, -1595, 7767, 3561, -6869, -5289, 5544, 6673, -3885, -7637, 1999, 8128, -8, -8131, -1972, 7653, 3819, -6735, -5435, 5437, 6727, -3844, -7636, 2047, 8115, -154, -8153, -1735, 7752, 3515, -6949, -5100, 5790, 6409, -4348, -7386, 2697, 7985, -928, -8191, -874, 8000, 2618, -7433, -4226, 6522, 5624, -5323, -6756, 3891, 7576, -2302, -8059, 624, 8187, 1064, -7970, -2695, 7421, 4198, -6575, -5520, 5471, 6608, -4163, -7431, 2703, 7958, -1156, -8183, -422, 8102, 1968, -7729, -3431, 7083, 4757, -6197, -5908, 5106, 6845, -3856, -7547, 2489, 7995, -1058, -8185, -395, 8115, 1819, -7798, -3174, 7249, 4420, -6494, -5526, 5558, 6461, -4478, -7207, 3284, 7748, -2016, -8077, 707, 8190, 604, -8095, -1887, 7798, 3107, -7315, -4240, 6662, 5258, -5864, -6145, 4941, 6882, -3921, -7461, 2826, 7872, -1688, -8116, 526, 8190, 629, -8103, -1759, 7859, 2839, -7473, -3854, 6953, 4784, -6318, -5619, 5580, 6345, -4760, -6958, 3872, 7447, -2936, -7815, 1967, 8056, -984, -8177, 0, 8176, 968, -8063, -1909, 7842, 2809, -7523, -3661, 7112, 4451, -6622, -5176, 6059, 5827, -5439, -6404, 4766, 6898, -4056, -7314, 3315, 7646, -2556, -7899, 1784, 8070, -1012, -8168, 243, 8189, 511, -8144, -1247, 8032, 1958, -7861, -2640, 7634, 3288, -7359, -3900, 7037, 4471, -6679, -5003, 6285, 5490, -5865, -5936, 5419, 6336, -4957, -6695, 4479, 7010, -3993, -7284, 3499, 7517, -3005, -7713, 2510, 7871, -2022, -7996, 1538, 8087, -1065, -8149, 601, 8182, -153, -8191, -283, 8176, 702, -8141, -1106, 8087, 1491, -8018, -1859, 7933, 2208, -7839, -2540, 7733, 2852, -7622, -3147, 7502, 3422, -7380, -3681, 7254, 3921, -7129, -4145, 7002, 4351, -6878, -4542, 6755, 4716, -6639, -4877, 6525, 5021, -6419, -5154, 6317, 5270, -6225, -5376, 6138, 5467, -6062, -5548, 5993, 5615, -5936, -5672, 5886, 5717, -5848, -5752, 5818, 5775, -5801, -5789, 5792, 5791, -5795, -5784, 5808, 5765, -5832, -5737, 5865, 5696, -5910, -5646, 5963, 5582, -6027, -5509, 6099, 5422, -6181, -5325, 6269, 5213, -6367, -5090, 6470, 4951, -6582, -4799, 6696, 4631, -6817, -4449, 6939, 4250, -7066, -4036, 7191, 3803, -7318, -3554, 7441, 3286, -7563, -3002, 7678, 2698, -7788, -2377, 7887, 2036, -7978, -1678, 8054, 1300, -8117, -907, 8160, 494, -8187, -68, 8189, -376, -8169, 831, 8121, -1301, -8046, 1778, 7937, -2266, -7797, 2757, 7620, -3253, -7406, 3746, 7152, -4237, -6858, 4719, 6521, -5191, -6142, 5644, 5718, -6079, -5252, 6485, 4742, -6863, -4191, 7203, 3598, -7503, -2969, 7753, 2302, -7954, -1606, 8095, 881, -8176, -136, 8187, -627, -8129, 1397, 7994, -2171, -7783, 2937, 7489, -3689, -7117, 4415, 6661, -5109, -6126, 5755, 5511, -6349, -4823, 6876, 4063, -7328, -3242, 7694, 2364, -7966, -1443, 8133, 486, -8191, 491, 8131, -1477, -7952, 2454, 7646, -3410, -7218, 4323, 6666, -5180, -5997, 5960, 5214, -6649, -4330, 7228, 3355, -7684, -2306, 8000, 1198, -8167, -54, 8174, -1108, -8016, 2260, 7687, -3381, -7193, 4441, 6532, -5417, -5720, 6280, 4764, -7009, -3686, 7578, 2506, -7971, -1252, 8168, -50, -8161, 1363, 7939, -2657, -7504, 3892, 6858, -5035, -6016, 6046, 4992, -6896, -3813, 7551, 2507, -7987, -1113, 8181, -331, -8123, 1778, 7803, -3184, -7228, 4498, 6404, -5675, -5357, 6667, 4113, -7438, -2714, 7950, 1202, -8181, 366, 8109, -1937, -7733, 3447, 7054, -4840, -6096, 6052, 4885, -7034, -3466, 7735, 1890, -8122, -223, 8167, -1470, -7861, 3112, 7207, -4632, -6227, 5955, 4954, -7018, -3444, 7761, 1758, -8145, 25, 8138, -1822, -7735, 3542, 6942, -5100, -5794, 6409, 4337, -7399, -2645, 8005, 797, -8190, 1106, 7930, -2965, -7234, 4671, 6125, -6129, -4662, 7245, 2918, -7951, -992, 8190, -1010, -7944, 2963, 7211, -4750, -6030, 6254, 4462, -7377, -2602, 8034, 559, -8177, 1533, 7782, -3539, -6867, 5320, 5480, -6753, -3710, 7727, 1669, -8170, 502, 8035, -2653, -7323, 4625, 6071, -6272, -4365, 7462, 2320, -8101, -87, 8123, -2168, -7520, 4267, 6323, -6046, -4618, 7351, 2531, -8072, -226, 8135, -2113, -7526, 4288, 6281, -6117, -4496, 7432, 2312, -8114, 85, 8087, -2490, -7345, 4685, 5938, -6473, -3985, 7677, 1653, -8181, 844, 7921, -3279, -6911, 5413, 5233, -7039, -3040, 7988, 534, -8156, 2036, 7511, -4418, -6107, 6364, 4071, -7669, -1606, 8185, -1042, -7848, 3592, 6675, -5775, -4783, 7346, 2360, -8126, 332, 8014, -3003, -7012, 5350, 5213, -7107, -2814, 8058, 78, -8085, 2680, 7166, -5139, -5399, 6999, 2978, -8032, -188, 8096, -2641, -7171, 5157, 5355, -7047, -2863, 8060, -5, -8059, 2883, 7025, -5407, -5079, 7238, 2458, -8130, 497, 7947, -3402, -6702, 5861, 4543, -7538, -1756, 8187, -1287, -7708, 4164, 6147, -6471, -3714, 7870, 739, -8150, 2354, 7253, -5121, -5295, 7149, 2548, -8130, 589, 7901, -3653, -6482, 6176, 4069, -7768, -1024, 8169, -2195, -7303, 5083, 5285, -7184, -2424, 8150, -839, -7814, 3978, 6210, -6486, -3586, 7938, 359, -8085, 2940, 6881, -5761, -4515, 7618, 1370, -8185, 2021, 7344, -5078, -5227, 7260, 2184, -8178, 1254, 7647, -4485, -5749, 6922, 2806, -8117, 658, 7834, -4016, -6109, 6644, 3243, -8046, 240, 7939, -3693, -6331, 6455, 3505, -7992, 4, 7988, -3528, -6430, 6373, 3600, -7974, -49, 7994, -3527, -6414, 6405, 3531, -7997, 80, 7959, -3689, -6284, 6548, 3296, -8054, 390, 7873, -4010, -6027, 6789, 2887, -8126, 882, 7714, -4476, -5626, 7104, 2296, -8182, 1550, 7450, -5067, -5055, 7460, 1513, -8179, 2382, 7040, -5749, -4287, 7805, 533, -8062, 3356, 6437, -6474, -3297, 8075, -637, -7764, 4430, 5594, -7174, -2070, 8190, -1970, -7217, 5540, 4469, -7760, -609, 8061, -3417, -6353, 6598, 3039, -8127, 1053, 7593, -4892, -5117, 7485, 1313, -8153, 2843, 6699, -6271, -3486, 8058, -659, -7719, 4640, 5319, -7395, -1485, 8164, -2764, -6723, 6273, 3441, -8076, 796, 7655, -4827, -5110, 7524, 1127, -8122, 3183, 6427, -6607, -2903, 8156, -1464, -7372, 5421, 4454, -7821, -234, 7945, -4068, -5740, 7183, 1830, -8181, 2633, 6739, -6324, -3272, 8119, -1195, -7460, 5311, 4523, -7815, -190, 7919, -4215, -5571, 7321, 1478, -8149, 3089, 6412, -6695, -2642, 8183, -1983, -7062, 5983, 3664, -8066, 927, 7535, -5230, -4544, 7831, 50, -7860, 4471, 5282, -7519, -936, 8059, -3737, -5890, 7160, 1718, -8162, 3048, 6377, -6784, -2398, 8190, -2423, -6763, 6413, 2971, -8171, 1872, 7058, -6068, -3445, 8120, -1405, -7280, 5763, 3822, -8059, 1023, 7440, -5512, -4111, 7996, -734, -7551, 5320, 4312, -7947, 535, 7618, -5197, -4434, 7915, -431, -7650, 5143, 4475, -7908, 417, 7647, -5163, -4440, 7923, -498, -7612, 5253, 4324, -7962, 670, 7538, -5414, -4128, 8016, -936, -7423, 5637, 3846, -8080, 1291, 7255, -5919, -3476, 8139, -1737, -7025) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L15_i
    );

    L15�31_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (5300, -4212, -8006, -921, 7416, 5663, -3801, -8089, -1351, 7231, 5943, -3463, -8138, -1686, 7074, 6148, -3202, -8164, -1927, 6955, 6285, -3025, -8176, -2077, 6883, 6360, -2933, -8181, -2137, 6859, 6375, -2927, -8180, -2107, 6886, 6332, -3008, -8174, -1986, 6963, 6228, -3175, -8159, -1775, 7084, 6060, -3425, -8127, -1471, 7243, 5821, -3754, -8070, -1073, 7430, 5503, -4156, -7975, -579, 7632, 5096, -4622, -7825, 10, 7832, 4591, -5140, -7604, 692, 8008, 3978, -5693, -7290, 1460, 8137, 3250, -6260, -6864, 2304, 8190, 2400, -6815, -6305, 3209, 8138, 1430, -7325, -5595, 4150, 7947, 346, -7754, -4721, 5095, 7586, -837, -8057, -3673, 6004, 7024, -2093, -8189, -2456, 6828, 6236, -3382, -8104, -1083, 7508, 5207, -4654, -7757, 414, 7983, 3935, -5844, -7111, 1988, 8187, 2437, -6874, -6141, 3571, 8059, 749, -7660, -4843, 5076, 7547, -1064, -8113, -3237, 6401, 6618, -2912, -8153, -1374, 7432, 5267, -4679, -7712, 659, 8055, 3525, -6228, -6751, 2739, 8164, 1465, -7412, -5271, 4711, 7681, -789, -8085, -3327, 6395, 6570, -3070, -8124, -1030, 7605, 4853, -5171, -7445, 1447, 8168, 2623, -6864, -6034, 3873, 7950, 54, -7926, -3956, 5982, 6890, -2610, -8167, -1375, 7498, 5019, -5064, -7473, 1451, 8173, 2485, -6980, -5836, 4185, 7836, -446, -8050, -3383, 6445, 6436, -3403, -8044, -387, 7862, 4076, -5954, -6861, 2752, 8143, 1033, -7665, -4584, 5546, 7143, -2258, -8182, -1495, 7498, 4921, -5255, -7314, 1932, 8190, 1774, -7391, -5106, 5093, 7393, -1782, -8191, -1875, 7356, 5145, -5075, -7393, 1808, 8190, 1796, -7403, -5042, 5197, 7311, -2013, -8188, -1541, 7521, 4790, -5456, -7140, 2390, 8164, 1101, -7696, -4380, 5834, 6854, -2934, -8095, -479, 7894, 3791, -6307, -6429, 3626, 7937, -330, -8076, -3010, 6834, 5823, -4443, -7646, 1315, 8183, 2017, -7365, -5004, 5340, 7160, -2457, -8149, -812, 7824, 3935, -6257, -6424, 3710, 7891, -595, -8127, -2600, 7107, 5381, -5008, -7333, 2159, 8169, 1000, -7785, -3999, 6249, 6393, -3806, -7846, 819, 8157, 2270, -7301, -5023, 5411, 7053, -2773, -8090, -242, 8000, 3207, -6815, -5723, 4709, 7451, -1981, -8176, -1000, 7813, 3833, -6427, -6154, 4211, 7666, -1466, -8191, -1455, 7674, 4176, -6198, -6364, 3957, 7754, -1243, -8189, -1611, 7629, 4255, -6160, -6380, 3965, 7740, -1318, -8191, -1470, 7692, 4074, -6318, -6203, 4234, 7621, -1689, -8185, -1031, 7843, 3623, -6650, -5810, 4745, 7361, -2347, -8125, -289, 8032, 2877, -7108, -5158, 5458, 6898, -3266, -7935, 757, 8173, 1811, -7607, -4190, 6300, 6147, -4397, -7507, 2083, 8147, 411, -8023, -2855, 7156, 5020, -5642, -6719, 3626, 7803, -1300, -8191, -1129, 7857, 3443, -6847, -5449, 5256, 6978, -3233, -7915, 950, 8187, 1395, -7790, -3614, 6764, 5527, -5207, -6992, 3247, 7899, -1049, -8191, -1218, 7855, 3376, -6932, -5269, 5497, 6760, -3671, -7750, 1589, 8175, 591, -8019, -2716, 7302, 4637, -6087, -6229, 4465, 7387, -2555, -8047, 488, 8171, 1595, -7767, -3563, 6868, 5289, -5544, -6674, 3884, 7636, -2000, -8129, 6, 8130, 1971, -7654, -3820, 6734, 5434, -5438, -6729, 3843, 7635, -2048, -8116, 153, 8152, 1734, -7753, -3516, 6948, 5100, -5791, -6410, 4346, 7385, -2697, -7987, 926, 8190, 874, -8001, -2619, 7431, 4225, -6523, -5625, 5321, 6756, -3892, -7577, 2301, 8058, -625, -8188, -1065, 7969, 2694, -7422, -4199, 6574, 5519, -5472, -6609, 4161, 7430, -2704, -7959, 1154, 8182, 422, -8103, -1970, 7728, 3430, -7083, -4758, 6196, 5907, -5107, -6846, 3854, 7547, -2490, -7996, 1056, 8184, 394, -8115, -1820, 7797, 3174, -7250, -4421, 6493, 5525, -5559, -6462, 4477, 7207, -3284, -7749, 2015, 8076, -707, -8191, -605, 8094, 1886, -7799, -3108, 7314, 4239, -6663, -5259, 5863, 6144, -4941, -6883, 3919, 7460, -2827, -7873, 1686, 8115, -527, -8191, -630, 8102, 1758, -7860, -2840, 7472, 3853, -6953, -4785, 6316, 5618, -5581, -6346, 4759, 6957, -3873, -7448, 2935, 7814, -1968, -8057, 983, 8176, -1, -8177, -969, 8062, 1909, -7843, -2810, 7522, 3660, -7112, -4452, 6621, 5175, -6060, -5828, 5438, 6403, -4767, -6899, 4055, 7313, -3316, -7647, 2555, 7898, -1785, -8071, 1011, 8167, -244, -8190, -512, 8143, 1247, -8032, -1959, 7860, 2640, -7635, -3289, 7358, 3899, -7038, -4472, 6678, 5002, -6286, -5491, 5864, 5935, -5420, -6337, 4956, 6694, -4480, -7011, 3992, 7284, -3500, -7518, 3004, 7712, -2511, -7872, 2020, 7995, -1539, -8088, 1064, 8148, -602, -8183, 152, 8190, 283, -8177, -703, 8140, 1105, -8088, -1492, 8017, 1859, -7934, -2209, 7838, 2539, -7734, -2853, 7621, 3146, -7503, -3423, 7379, 3680, -7255, -3922, 7128, 4144, -7003, -4352, 6877, 4541, -6756, -4717, 6638, 4876, -6526, -5022, 6418, 5153, -6318, -5271, 6224, 5375, -6139, -5468, 6061, 5547, -5994, -5616, 5935, 5672, -5887, -5718, 5847, 5751, -5819, -5776, 5800, 5788, -5793, -5792, 5794, 5783, -5809, -5766, 5831, 5736, -5866, -5697, 5909, 5645, -5964, -5583, 6026, 5508, -6100, -5423, 6180, 5324, -6270, -5214, 6366, 5089, -6471, -4952, 6581, 4798, -6697, -4632, 6816, 4448, -6940, -4250, 7065, 4034, -7192, -3804, 7317, 3553, -7442, -3287, 7562, 3001, -7679, -2699, 7787, 2376, -7888, -2036, 7977, 1677, -8055, -1301, 8116, 906, -8161, -495, 8186, 67, -8190, 375, 8168, -832, -8122, 1300, 8045, -1779, -7938, 2265, 7796, -2758, -7620, 3252, 7405, -3747, -7153, 4236, 6857, -4720, -6522, 5190, 6141, -5645, -5719, 6078, 5251, -6487, -4743, 6862, 4190, -7204, -3599, 7502, 2968, -7754, -2303, 7953, 1605, -8096, -882, 8175, 135, -8188, 626, 8128, -1398, -7995, 2170, 7782, -2938, -7490, 3688, 7116, -4416, -6662, 5108, 6125, -5756, -5511, 6348, 4821, -6877, -4064, 7327, 3241, -7695, -2365, 7965, 1442, -8134, -487, 8190, -492, -8132, 1476, 7951, -2455, -7647, 3409, 7217, -4324, -6667, 5179, 5995, -5961, -5215, 6648, 4329, -7229, -3356, 7683, 2305, -8001, -1199, 8166, 52, -8175, 1108, 8015, -2262, -7688, 3380, 7191, -4442, -6533, 5416, 5718, -6281, -4764, 7008, 3685, -7579, -2507, 7970, 1251, -8169, 49, 8160, -1365, -7940, 2657, 7503, -3893, -6859, 5034, 6015, -6047, -4993, 6895, 3812, -7552, -2508, 7986, 1112, -8182, 331, 8122, -1779, -7804, 3184, 7226, -4499, -6405, 5674, 5356, -6668, -4114, 7438, 2713, -7951, -1203, 8180, -367, -8110, 1936, 7731, -3449, -7055, 4839, 6095, -6053, -4885, 7033, 3465, -7736, -1891, 8121, 222, -8168, 1469, 7860, -3113, -7208, 4631, 6226, -5956, -4955, 7017, 3443, -7762, -1758, 8144, -26, -8139, 1821, 7734, -3543, -6943, 5100, 5792, -6411, -4338, 7398, 2643, -8006, -797, 8189, -1107, -7931, 2964, 7233, -4673, -6126, 6129, 4661, -7247, -2918, 7950, 990, -8191, 1009, 7943, -2964, -7211, 4750, 6029, -6255, -4462, 7376, 2600, -8035, -559, 8176, -1534, -7783, 3538, 6866, -5321, -5481, 6752, 3709, -7729, -1669, 8169, -503, -8036, 2653, 7322, -4626, -6072, 6272, 4364, -7464, -2320, 8100, 86, -8124, 2168, 7519, -4269, -6323, 6045, 4617, -7352, -2531, 8071, 225, -8136, 2113, 7525, -4290, -6281, 6116, 4494, -7433, -2312, 8113, -86, -8088, 2490, 7344, -4687, -5938, 6472, 3983, -7679, -1653, 8180, -846, -7922, 3278, 6910, -5414, -5233, 7039, 3038, -7989, -535, 8155, -2037, -7512, 4418, 6106, -6365, -4071, 7669, 1604, -8186, 1042, 7847, -3594, -6676, 5775, 4781, -7347, -2361, 8126, -333, -8015, 3003, 7010, -5352, -5214, 7106, 2813, -8059, -78, 8084, -2681, -7167, 5138, 5398, -7000, -2979, 8031, 187, -8096, 2640, 7170, -5158, -5355, 7046, 2861, -8062, 4, 8058, -2885, -7025, 5406, 5077, -7239, -2459, 8129, -498, -7948, 3401, 6701, -5862, -4544, 7537, 1755, -8188, 1287, 7707, -4166, -6148, 6471, 3713, -7871, -739, 8149, -2356, -7253, 5121, 5294, -7150, -2548, 8129, -590, -7901, 3652, 6480, -6177, -4070, 7767, 1022, -8170, 2195, 7301, -5085, -5286, 7184, 2422, -8151, 839, 7813, -3980, -6210, 6485, 3585, -7940, -359, 8084, -2941, -6881, 5761, 4513, -7619, -1370, 8184, -2022, -7344, 5077, 5225, -7262, -2185, 8177, -1256, -7648, 4485, 5748, -6923, -2806, 8116, -660, -7835, 4016, 6108, -6645, -3243, 8045, -242, -7940, 3693, 6329, -6457, -3505, 7991, -6, -7989, 3528, 6428, -6375, -3600, 7974, 47, -7995, 3527, 6413, -6407, -3531, 7996, -81, -7960, 3689, 6282, -6549, -3296, 8053, -392, -7874, 4010, 6025, -6790, -2887, 8125, -884, -7715, 4476, 5624, -7106, -2296, 8181, -1552, -7451, 5067, 5053, -7461, -1513, 8178, -2384, -7041, 5749, 4285, -7806, -533, 8061, -3358, -6438, 6474, 3295, -8076, 636, 7763, -4431, -5594, 7173, 2068, -8191, 1970, 7216, -5542, -4469, 7759, 607, -8062, 3417, 6351, -6600, -3039, 8126, -1055, -7594, 4891, 5115, -7486, -1313, 8152, -2845, -6700, 6270, 3485, -8060, 659, 7718, -4642, -5319, 7394, 1483, -8165, 2764, 6722, -6274, -3441, 8075, -798, -7656, 4827, 5108, -7526, -1127, 8121, -3185, -6428, 6607, 2901, -8157, 1464, 7370, -5423, -4454, 7820, 232, -7946, 4068, 5738, -7185, -1830, 8180, -2635, -6740, 6323, 3270, -8120, 1195, 7459, -5313, -4523, 7814, 188, -7919, 4215, 5569, -7323, -1478, 8147, -3091, -6412, 6695, 2640, -8184, 1983, 7060, -5984, -3664, 8065, -929, -7536, 5230, 4542, -7832, -50, 7859, -4473, -5282, 7519, 934, -8060, 3737, 5888, -7161, -1718, 8161, -3050, -6377, 6784, 2395, -8191, 2423, 6761, -6414, -2971, 8170, -1874, -7058, 6068, 3443, -8121, 1405, 7279, -5765, -3822, 8058, -1025, -7440, 5512, 4109, -7997, 735, 7549, -5322, -4312, 7947, -537, -7618, 5197, 4432, -7917, 431, 7649, -5145, -4475, 7908, -419, -7648, 5163, 4438, -7924, 499, 7611, -5255, -4324, 7961, -673, -7539, 5413, 4126, -8017, 937, 7422, -5639, -3846, 8079, -1294, -7255, 5918, 3474, -8140, 1737, 7024) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L15�31_i
    );

    L15�32_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-5300, 4212, 8004, 919, -7418, -5663, 3801, 8088, 1349, -7232, -5943, 3463, 8137, 1683, -7075, -6148, 3202, 8163, 1925, -6957, -6285, 3025, 8175, 2075, -6884, -6360, 2933, 8180, 2135, -6861, -6375, 2927, 8179, 2105, -6888, -6332, 3008, 8173, 1984, -6964, -6228, 3175, 8158, 1773, -7085, -6060, 3425, 8126, 1469, -7245, -5821, 3754, 8069, 1070, -7432, -5503, 4156, 7974, 577, -7634, -5096, 4622, 7824, -12, -7833, -4591, 5139, 7602, -694, -8009, -3978, 5693, 7289, -1462, -8138, -3250, 6260, 6862, -2306, -8191, -2400, 6815, 6304, -3211, -8139, -1430, 7325, 5594, -4152, -7948, -346, 7753, 4719, -5097, -7586, 837, 8056, 3672, -6006, -7024, 2093, 8188, 2454, -6829, -6236, 3382, 8103, 1081, -7510, -5207, 4654, 7756, -416, -7984, -3935, 5844, 7109, -1990, -8188, -2437, 6874, 6140, -3573, -8060, -749, 7659, 4841, -5078, -7547, 1064, 8113, 3235, -6402, -6618, 2912, 8152, 1372, -7433, -5267, 4679, 7710, -661, -8056, -3525, 6228, 6749, -2741, -8165, -1465, 7412, 5270, -4713, -7682, 789, 8085, 3325, -6397, -6571, 3070, 8122, 1028, -7607, -4853, 5171, 7444, -1449, -8169, -2623, 6864, 6032, -3875, -7951, -54, 7925, 3954, -5984, -6890, 2610, 8166, 1373, -7499, -5019, 5064, 7471, -1453, -8174, -2485, 6980, 5834, -4186, -7837, 445, 8050, 3381, -6446, -6436, 3403, 8042, 385, -7863, -4076, 5954, 6860, -2754, -8144, -1033, 7665, 4582, -5548, -7143, 2258, 8181, 1494, -7499, -4921, 5254, 7313, -1933, -8191, -1774, 7390, 5104, -5095, -7394, 1782, 8190, 1873, -7358, -5145, 5075, 7392, -1810, -8191, -1796, 7402, 5041, -5199, -7312, 2013, 8187, 1539, -7522, -4791, 5456, 7139, -2391, -8165, -1102, 7695, 4379, -5835, -6855, 2933, 8094, 477, -7895, -3792, 6307, 6427, -3627, -7938, 330, 8075, 3008, -6835, -5824, 4443, 7645, -1317, -8184, -2017, 7364, 5003, -5341, -7160, 2456, 8147, 810, -7825, -3935, 6257, 6422, -3711, -7892, 595, 8126, 2598, -7109, -5381, 5008, 7331, -2160, -8170, -1001, 7784, 3997, -6250, -6393, 3805, 7845, -821, -8158, -2270, 7300, 5021, -5413, -7054, 2772, 8089, 240, -8001, -3207, 6815, 5721, -4710, -7452, 1980, 8175, 999, -7814, -3834, 6426, 6153, -4212, -7667, 1465, 8190, 1453, -7675, -4177, 6197, 6363, -3959, -7754, 1243, 8188, 1609, -7631, -4255, 6159, 6378, -3967, -7741, 1318, 8190, 1469, -7693, -4074, 6317, 6201, -4235, -7621, 1689, 8184, 1030, -7844, -3623, 6649, 5808, -4747, -7361, 2346, 8124, 287, -8033, -2878, 7107, 5156, -5460, -6898, 3266, 7933, -759, -8174, -1812, 7606, 4188, -6302, -6148, 4396, 7506, -2085, -8148, -411, 8022, 2853, -7157, -5021, 5641, 6718, -3627, -7804, 1300, 8190, 1127, -7858, -3443, 6847, 5448, -5258, -6979, 3233, 7913, -952, -8188, -1395, 7790, 3612, -6766, -5528, 5206, 6991, -3249, -7899, 1048, 8190, 1216, -7856, -3376, 6931, 5268, -5498, -6761, 3670, 7749, -1591, -8176, -591, 8019, 2715, -7303, -4637, 6087, 6227, -4466, -7388, 2555, 8046, -490, -8172, -1595, 7767, 3561, -6869, -5289, 5544, 6673, -3885, -7637, 1999, 8128, -8, -8131, -1972, 7653, 3819, -6735, -5435, 5437, 6727, -3844, -7636, 2047, 8115, -154, -8153, -1735, 7752, 3515, -6949, -5100, 5790, 6409, -4348, -7386, 2697, 7985, -928, -8191, -874, 8000, 2618, -7433, -4226, 6522, 5624, -5323, -6756, 3891, 7576, -2302, -8059, 624, 8187, 1064, -7970, -2695, 7421, 4198, -6575, -5520, 5471, 6608, -4163, -7431, 2703, 7958, -1156, -8183, -422, 8102, 1968, -7729, -3431, 7083, 4757, -6197, -5908, 5106, 6845, -3856, -7547, 2489, 7995, -1058, -8185, -395, 8115, 1819, -7798, -3174, 7249, 4420, -6494, -5526, 5558, 6461, -4478, -7207, 3284, 7748, -2016, -8077, 707, 8190, 604, -8095, -1887, 7798, 3107, -7315, -4240, 6662, 5258, -5864, -6145, 4941, 6882, -3921, -7461, 2826, 7872, -1688, -8116, 526, 8190, 629, -8103, -1759, 7859, 2839, -7473, -3854, 6953, 4784, -6318, -5619, 5580, 6345, -4760, -6958, 3872, 7447, -2936, -7815, 1967, 8056, -984, -8177, 0, 8176, 968, -8063, -1909, 7842, 2809, -7523, -3661, 7112, 4451, -6622, -5176, 6059, 5827, -5439, -6404, 4766, 6898, -4056, -7314, 3315, 7646, -2556, -7899, 1784, 8070, -1012, -8168, 243, 8189, 511, -8144, -1247, 8032, 1958, -7861, -2640, 7634, 3288, -7359, -3900, 7037, 4471, -6679, -5003, 6285, 5490, -5865, -5936, 5419, 6336, -4957, -6695, 4479, 7010, -3993, -7284, 3499, 7517, -3005, -7713, 2510, 7871, -2022, -7996, 1538, 8087, -1065, -8149, 601, 8182, -153, -8191, -283, 8176, 702, -8141, -1106, 8087, 1491, -8018, -1859, 7933, 2208, -7839, -2540, 7733, 2852, -7622, -3147, 7502, 3422, -7380, -3681, 7254, 3921, -7129, -4145, 7002, 4351, -6878, -4542, 6755, 4716, -6639, -4877, 6525, 5021, -6419, -5154, 6317, 5270, -6225, -5376, 6138, 5467, -6062, -5548, 5993, 5615, -5936, -5672, 5886, 5717, -5848, -5752, 5818, 5775, -5801, -5789, 5792, 5791, -5795, -5784, 5808, 5765, -5832, -5737, 5865, 5696, -5910, -5646, 5963, 5582, -6027, -5509, 6099, 5422, -6181, -5325, 6269, 5213, -6367, -5090, 6470, 4951, -6582, -4799, 6696, 4631, -6817, -4449, 6939, 4250, -7066, -4036, 7191, 3803, -7318, -3554, 7441, 3286, -7563, -3002, 7678, 2698, -7788, -2377, 7887, 2036, -7978, -1678, 8054, 1300, -8117, -907, 8160, 494, -8187, -68, 8189, -376, -8169, 831, 8121, -1301, -8046, 1778, 7937, -2266, -7797, 2757, 7620, -3253, -7406, 3746, 7152, -4237, -6858, 4719, 6521, -5191, -6142, 5644, 5718, -6079, -5252, 6485, 4742, -6863, -4191, 7203, 3598, -7503, -2969, 7753, 2302, -7954, -1606, 8095, 881, -8176, -136, 8187, -627, -8129, 1397, 7994, -2171, -7783, 2937, 7489, -3689, -7117, 4415, 6661, -5109, -6126, 5755, 5511, -6349, -4823, 6876, 4063, -7328, -3242, 7694, 2364, -7966, -1443, 8133, 486, -8191, 491, 8131, -1477, -7952, 2454, 7646, -3410, -7218, 4323, 6666, -5180, -5997, 5960, 5214, -6649, -4330, 7228, 3355, -7684, -2306, 8000, 1198, -8167, -54, 8174, -1108, -8016, 2260, 7687, -3381, -7193, 4441, 6532, -5417, -5720, 6280, 4764, -7009, -3686, 7578, 2506, -7971, -1252, 8168, -50, -8161, 1363, 7939, -2657, -7504, 3892, 6858, -5035, -6016, 6046, 4992, -6896, -3813, 7551, 2507, -7987, -1113, 8181, -331, -8123, 1778, 7803, -3184, -7228, 4498, 6404, -5675, -5357, 6667, 4113, -7438, -2714, 7950, 1202, -8181, 366, 8109, -1937, -7733, 3447, 7054, -4840, -6096, 6052, 4885, -7034, -3466, 7735, 1890, -8122, -223, 8167, -1470, -7861, 3112, 7207, -4632, -6227, 5955, 4954, -7018, -3444, 7761, 1758, -8145, 25, 8138, -1822, -7735, 3542, 6942, -5100, -5794, 6409, 4337, -7399, -2645, 8005, 797, -8190, 1106, 7930, -2965, -7234, 4671, 6125, -6129, -4662, 7245, 2918, -7951, -992, 8190, -1010, -7944, 2963, 7211, -4750, -6030, 6254, 4462, -7377, -2602, 8034, 559, -8177, 1533, 7782, -3539, -6867, 5320, 5480, -6753, -3710, 7727, 1669, -8170, 502, 8035, -2653, -7323, 4625, 6071, -6272, -4365, 7462, 2320, -8101, -87, 8123, -2168, -7520, 4267, 6323, -6046, -4618, 7351, 2531, -8072, -226, 8135, -2113, -7526, 4288, 6281, -6117, -4496, 7432, 2312, -8114, 85, 8087, -2490, -7345, 4685, 5938, -6473, -3985, 7677, 1653, -8181, 844, 7921, -3279, -6911, 5413, 5233, -7039, -3040, 7988, 534, -8156, 2036, 7511, -4418, -6107, 6364, 4071, -7669, -1606, 8185, -1042, -7848, 3592, 6675, -5775, -4783, 7346, 2360, -8126, 332, 8014, -3003, -7012, 5350, 5213, -7107, -2814, 8058, 78, -8085, 2680, 7166, -5139, -5399, 6999, 2978, -8032, -188, 8096, -2641, -7171, 5157, 5355, -7047, -2863, 8060, -5, -8059, 2883, 7025, -5407, -5079, 7238, 2458, -8130, 497, 7947, -3402, -6702, 5861, 4543, -7538, -1756, 8187, -1287, -7708, 4164, 6147, -6471, -3714, 7870, 739, -8150, 2354, 7253, -5121, -5295, 7149, 2548, -8130, 589, 7901, -3653, -6482, 6176, 4069, -7768, -1024, 8169, -2195, -7303, 5083, 5285, -7184, -2424, 8150, -839, -7814, 3978, 6210, -6486, -3586, 7938, 359, -8085, 2940, 6881, -5761, -4515, 7618, 1370, -8185, 2021, 7344, -5078, -5227, 7260, 2184, -8178, 1254, 7647, -4485, -5749, 6922, 2806, -8117, 658, 7834, -4016, -6109, 6644, 3243, -8046, 240, 7939, -3693, -6331, 6455, 3505, -7992, 4, 7988, -3528, -6430, 6373, 3600, -7974, -49, 7994, -3527, -6414, 6405, 3531, -7997, 80, 7959, -3689, -6284, 6548, 3296, -8054, 390, 7873, -4010, -6027, 6789, 2887, -8126, 882, 7714, -4476, -5626, 7104, 2296, -8182, 1550, 7450, -5067, -5055, 7460, 1513, -8179, 2382, 7040, -5749, -4287, 7805, 533, -8062, 3356, 6437, -6474, -3297, 8075, -637, -7764, 4430, 5594, -7174, -2070, 8190, -1970, -7217, 5540, 4469, -7760, -609, 8061, -3417, -6353, 6598, 3039, -8127, 1053, 7593, -4892, -5117, 7485, 1313, -8153, 2843, 6699, -6271, -3486, 8058, -659, -7719, 4640, 5319, -7395, -1485, 8164, -2764, -6723, 6273, 3441, -8076, 796, 7655, -4827, -5110, 7524, 1127, -8122, 3183, 6427, -6607, -2903, 8156, -1464, -7372, 5421, 4454, -7821, -234, 7945, -4068, -5740, 7183, 1830, -8181, 2633, 6739, -6324, -3272, 8119, -1195, -7460, 5311, 4523, -7815, -190, 7919, -4215, -5571, 7321, 1478, -8149, 3089, 6412, -6695, -2642, 8183, -1983, -7062, 5983, 3664, -8066, 927, 7535, -5230, -4544, 7831, 50, -7860, 4471, 5282, -7519, -936, 8059, -3737, -5890, 7160, 1718, -8162, 3048, 6377, -6784, -2398, 8190, -2423, -6763, 6413, 2971, -8171, 1872, 7058, -6068, -3445, 8120, -1405, -7280, 5763, 3822, -8059, 1023, 7440, -5512, -4111, 7996, -734, -7551, 5320, 4312, -7947, 535, 7618, -5197, -4434, 7915, -431, -7650, 5143, 4475, -7908, 417, 7647, -5163, -4440, 7923, -498, -7612, 5253, 4324, -7962, 670, 7538, -5414, -4128, 8016, -936, -7423, 5637, 3846, -8080, 1291, 7255, -5919, -3476, 8139, -1737, -7025) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L15�32_i
    );

    L15�33_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (5300, -4212, -8006, -921, 7416, 5663, -3801, -8089, -1351, 7231, 5943, -3463, -8138, -1686, 7074, 6148, -3202, -8164, -1927, 6955, 6285, -3025, -8176, -2077, 6883, 6360, -2933, -8181, -2137, 6859, 6375, -2927, -8180, -2107, 6886, 6332, -3008, -8174, -1986, 6963, 6228, -3175, -8159, -1775, 7084, 6060, -3425, -8127, -1471, 7243, 5821, -3754, -8070, -1073, 7430, 5503, -4156, -7975, -579, 7632, 5096, -4622, -7825, 10, 7832, 4591, -5140, -7604, 692, 8008, 3978, -5693, -7290, 1460, 8137, 3250, -6260, -6864, 2304, 8190, 2400, -6815, -6305, 3209, 8138, 1430, -7325, -5595, 4150, 7947, 346, -7754, -4721, 5095, 7586, -837, -8057, -3673, 6004, 7024, -2093, -8189, -2456, 6828, 6236, -3382, -8104, -1083, 7508, 5207, -4654, -7757, 414, 7983, 3935, -5844, -7111, 1988, 8187, 2437, -6874, -6141, 3571, 8059, 749, -7660, -4843, 5076, 7547, -1064, -8113, -3237, 6401, 6618, -2912, -8153, -1374, 7432, 5267, -4679, -7712, 659, 8055, 3525, -6228, -6751, 2739, 8164, 1465, -7412, -5271, 4711, 7681, -789, -8085, -3327, 6395, 6570, -3070, -8124, -1030, 7605, 4853, -5171, -7445, 1447, 8168, 2623, -6864, -6034, 3873, 7950, 54, -7926, -3956, 5982, 6890, -2610, -8167, -1375, 7498, 5019, -5064, -7473, 1451, 8173, 2485, -6980, -5836, 4185, 7836, -446, -8050, -3383, 6445, 6436, -3403, -8044, -387, 7862, 4076, -5954, -6861, 2752, 8143, 1033, -7665, -4584, 5546, 7143, -2258, -8182, -1495, 7498, 4921, -5255, -7314, 1932, 8190, 1774, -7391, -5106, 5093, 7393, -1782, -8191, -1875, 7356, 5145, -5075, -7393, 1808, 8190, 1796, -7403, -5042, 5197, 7311, -2013, -8188, -1541, 7521, 4790, -5456, -7140, 2390, 8164, 1101, -7696, -4380, 5834, 6854, -2934, -8095, -479, 7894, 3791, -6307, -6429, 3626, 7937, -330, -8076, -3010, 6834, 5823, -4443, -7646, 1315, 8183, 2017, -7365, -5004, 5340, 7160, -2457, -8149, -812, 7824, 3935, -6257, -6424, 3710, 7891, -595, -8127, -2600, 7107, 5381, -5008, -7333, 2159, 8169, 1000, -7785, -3999, 6249, 6393, -3806, -7846, 819, 8157, 2270, -7301, -5023, 5411, 7053, -2773, -8090, -242, 8000, 3207, -6815, -5723, 4709, 7451, -1981, -8176, -1000, 7813, 3833, -6427, -6154, 4211, 7666, -1466, -8191, -1455, 7674, 4176, -6198, -6364, 3957, 7754, -1243, -8189, -1611, 7629, 4255, -6160, -6380, 3965, 7740, -1318, -8191, -1470, 7692, 4074, -6318, -6203, 4234, 7621, -1689, -8185, -1031, 7843, 3623, -6650, -5810, 4745, 7361, -2347, -8125, -289, 8032, 2877, -7108, -5158, 5458, 6898, -3266, -7935, 757, 8173, 1811, -7607, -4190, 6300, 6147, -4397, -7507, 2083, 8147, 411, -8023, -2855, 7156, 5020, -5642, -6719, 3626, 7803, -1300, -8191, -1129, 7857, 3443, -6847, -5449, 5256, 6978, -3233, -7915, 950, 8187, 1395, -7790, -3614, 6764, 5527, -5207, -6992, 3247, 7899, -1049, -8191, -1218, 7855, 3376, -6932, -5269, 5497, 6760, -3671, -7750, 1589, 8175, 591, -8019, -2716, 7302, 4637, -6087, -6229, 4465, 7387, -2555, -8047, 488, 8171, 1595, -7767, -3563, 6868, 5289, -5544, -6674, 3884, 7636, -2000, -8129, 6, 8130, 1971, -7654, -3820, 6734, 5434, -5438, -6729, 3843, 7635, -2048, -8116, 153, 8152, 1734, -7753, -3516, 6948, 5100, -5791, -6410, 4346, 7385, -2697, -7987, 926, 8190, 874, -8001, -2619, 7431, 4225, -6523, -5625, 5321, 6756, -3892, -7577, 2301, 8058, -625, -8188, -1065, 7969, 2694, -7422, -4199, 6574, 5519, -5472, -6609, 4161, 7430, -2704, -7959, 1154, 8182, 422, -8103, -1970, 7728, 3430, -7083, -4758, 6196, 5907, -5107, -6846, 3854, 7547, -2490, -7996, 1056, 8184, 394, -8115, -1820, 7797, 3174, -7250, -4421, 6493, 5525, -5559, -6462, 4477, 7207, -3284, -7749, 2015, 8076, -707, -8191, -605, 8094, 1886, -7799, -3108, 7314, 4239, -6663, -5259, 5863, 6144, -4941, -6883, 3919, 7460, -2827, -7873, 1686, 8115, -527, -8191, -630, 8102, 1758, -7860, -2840, 7472, 3853, -6953, -4785, 6316, 5618, -5581, -6346, 4759, 6957, -3873, -7448, 2935, 7814, -1968, -8057, 983, 8176, -1, -8177, -969, 8062, 1909, -7843, -2810, 7522, 3660, -7112, -4452, 6621, 5175, -6060, -5828, 5438, 6403, -4767, -6899, 4055, 7313, -3316, -7647, 2555, 7898, -1785, -8071, 1011, 8167, -244, -8190, -512, 8143, 1247, -8032, -1959, 7860, 2640, -7635, -3289, 7358, 3899, -7038, -4472, 6678, 5002, -6286, -5491, 5864, 5935, -5420, -6337, 4956, 6694, -4480, -7011, 3992, 7284, -3500, -7518, 3004, 7712, -2511, -7872, 2020, 7995, -1539, -8088, 1064, 8148, -602, -8183, 152, 8190, 283, -8177, -703, 8140, 1105, -8088, -1492, 8017, 1859, -7934, -2209, 7838, 2539, -7734, -2853, 7621, 3146, -7503, -3423, 7379, 3680, -7255, -3922, 7128, 4144, -7003, -4352, 6877, 4541, -6756, -4717, 6638, 4876, -6526, -5022, 6418, 5153, -6318, -5271, 6224, 5375, -6139, -5468, 6061, 5547, -5994, -5616, 5935, 5672, -5887, -5718, 5847, 5751, -5819, -5776, 5800, 5788, -5793, -5792, 5794, 5783, -5809, -5766, 5831, 5736, -5866, -5697, 5909, 5645, -5964, -5583, 6026, 5508, -6100, -5423, 6180, 5324, -6270, -5214, 6366, 5089, -6471, -4952, 6581, 4798, -6697, -4632, 6816, 4448, -6940, -4250, 7065, 4034, -7192, -3804, 7317, 3553, -7442, -3287, 7562, 3001, -7679, -2699, 7787, 2376, -7888, -2036, 7977, 1677, -8055, -1301, 8116, 906, -8161, -495, 8186, 67, -8190, 375, 8168, -832, -8122, 1300, 8045, -1779, -7938, 2265, 7796, -2758, -7620, 3252, 7405, -3747, -7153, 4236, 6857, -4720, -6522, 5190, 6141, -5645, -5719, 6078, 5251, -6487, -4743, 6862, 4190, -7204, -3599, 7502, 2968, -7754, -2303, 7953, 1605, -8096, -882, 8175, 135, -8188, 626, 8128, -1398, -7995, 2170, 7782, -2938, -7490, 3688, 7116, -4416, -6662, 5108, 6125, -5756, -5511, 6348, 4821, -6877, -4064, 7327, 3241, -7695, -2365, 7965, 1442, -8134, -487, 8190, -492, -8132, 1476, 7951, -2455, -7647, 3409, 7217, -4324, -6667, 5179, 5995, -5961, -5215, 6648, 4329, -7229, -3356, 7683, 2305, -8001, -1199, 8166, 52, -8175, 1108, 8015, -2262, -7688, 3380, 7191, -4442, -6533, 5416, 5718, -6281, -4764, 7008, 3685, -7579, -2507, 7970, 1251, -8169, 49, 8160, -1365, -7940, 2657, 7503, -3893, -6859, 5034, 6015, -6047, -4993, 6895, 3812, -7552, -2508, 7986, 1112, -8182, 331, 8122, -1779, -7804, 3184, 7226, -4499, -6405, 5674, 5356, -6668, -4114, 7438, 2713, -7951, -1203, 8180, -367, -8110, 1936, 7731, -3449, -7055, 4839, 6095, -6053, -4885, 7033, 3465, -7736, -1891, 8121, 222, -8168, 1469, 7860, -3113, -7208, 4631, 6226, -5956, -4955, 7017, 3443, -7762, -1758, 8144, -26, -8139, 1821, 7734, -3543, -6943, 5100, 5792, -6411, -4338, 7398, 2643, -8006, -797, 8189, -1107, -7931, 2964, 7233, -4673, -6126, 6129, 4661, -7247, -2918, 7950, 990, -8191, 1009, 7943, -2964, -7211, 4750, 6029, -6255, -4462, 7376, 2600, -8035, -559, 8176, -1534, -7783, 3538, 6866, -5321, -5481, 6752, 3709, -7729, -1669, 8169, -503, -8036, 2653, 7322, -4626, -6072, 6272, 4364, -7464, -2320, 8100, 86, -8124, 2168, 7519, -4269, -6323, 6045, 4617, -7352, -2531, 8071, 225, -8136, 2113, 7525, -4290, -6281, 6116, 4494, -7433, -2312, 8113, -86, -8088, 2490, 7344, -4687, -5938, 6472, 3983, -7679, -1653, 8180, -846, -7922, 3278, 6910, -5414, -5233, 7039, 3038, -7989, -535, 8155, -2037, -7512, 4418, 6106, -6365, -4071, 7669, 1604, -8186, 1042, 7847, -3594, -6676, 5775, 4781, -7347, -2361, 8126, -333, -8015, 3003, 7010, -5352, -5214, 7106, 2813, -8059, -78, 8084, -2681, -7167, 5138, 5398, -7000, -2979, 8031, 187, -8096, 2640, 7170, -5158, -5355, 7046, 2861, -8062, 4, 8058, -2885, -7025, 5406, 5077, -7239, -2459, 8129, -498, -7948, 3401, 6701, -5862, -4544, 7537, 1755, -8188, 1287, 7707, -4166, -6148, 6471, 3713, -7871, -739, 8149, -2356, -7253, 5121, 5294, -7150, -2548, 8129, -590, -7901, 3652, 6480, -6177, -4070, 7767, 1022, -8170, 2195, 7301, -5085, -5286, 7184, 2422, -8151, 839, 7813, -3980, -6210, 6485, 3585, -7940, -359, 8084, -2941, -6881, 5761, 4513, -7619, -1370, 8184, -2022, -7344, 5077, 5225, -7262, -2185, 8177, -1256, -7648, 4485, 5748, -6923, -2806, 8116, -660, -7835, 4016, 6108, -6645, -3243, 8045, -242, -7940, 3693, 6329, -6457, -3505, 7991, -6, -7989, 3528, 6428, -6375, -3600, 7974, 47, -7995, 3527, 6413, -6407, -3531, 7996, -81, -7960, 3689, 6282, -6549, -3296, 8053, -392, -7874, 4010, 6025, -6790, -2887, 8125, -884, -7715, 4476, 5624, -7106, -2296, 8181, -1552, -7451, 5067, 5053, -7461, -1513, 8178, -2384, -7041, 5749, 4285, -7806, -533, 8061, -3358, -6438, 6474, 3295, -8076, 636, 7763, -4431, -5594, 7173, 2068, -8191, 1970, 7216, -5542, -4469, 7759, 607, -8062, 3417, 6351, -6600, -3039, 8126, -1055, -7594, 4891, 5115, -7486, -1313, 8152, -2845, -6700, 6270, 3485, -8060, 659, 7718, -4642, -5319, 7394, 1483, -8165, 2764, 6722, -6274, -3441, 8075, -798, -7656, 4827, 5108, -7526, -1127, 8121, -3185, -6428, 6607, 2901, -8157, 1464, 7370, -5423, -4454, 7820, 232, -7946, 4068, 5738, -7185, -1830, 8180, -2635, -6740, 6323, 3270, -8120, 1195, 7459, -5313, -4523, 7814, 188, -7919, 4215, 5569, -7323, -1478, 8147, -3091, -6412, 6695, 2640, -8184, 1983, 7060, -5984, -3664, 8065, -929, -7536, 5230, 4542, -7832, -50, 7859, -4473, -5282, 7519, 934, -8060, 3737, 5888, -7161, -1718, 8161, -3050, -6377, 6784, 2395, -8191, 2423, 6761, -6414, -2971, 8170, -1874, -7058, 6068, 3443, -8121, 1405, 7279, -5765, -3822, 8058, -1025, -7440, 5512, 4109, -7997, 735, 7549, -5322, -4312, 7947, -537, -7618, 5197, 4432, -7917, 431, 7649, -5145, -4475, 7908, -419, -7648, 5163, 4438, -7924, 499, 7611, -5255, -4324, 7961, -673, -7539, 5413, 4126, -8017, 937, 7422, -5639, -3846, 8079, -1294, -7255, 5918, 3474, -8140, 1737, 7024) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L15�33_i
    );

    L21_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (5500, 7514, -675, -7949, -4422, 5117, 7696, -198, -7824, -4795, 4767, 7831, 215, -7696, -5104, 4457, 7929, 564, -7574, -5352, 4194, 7999, 846, -7467, -5545, 3982, 8045, 1064, -7380, -5686, 3823, 8075, 1217, -7317, -5778, 3720, 8092, 1306, -7282, -5823, 3675, 8098, 1331, -7277, -5823, 3687, 8093, 1292, -7300, -5777, 3756, 8079, 1190, -7353, -5684, 3883, 8052, 1023, -7431, -5542, 4064, 8009, 791, -7531, -5349, 4298, 7944, 494, -7648, -5100, 4581, 7852, 132, -7774, -4790, 4908, 7724, -296, -7902, -4415, 5273, 7552, -786, -8020, -3971, 5667, 7325, -1338, -8116, -3452, 6082, 7032, -1946, -8178, -2855, 6504, 6664, -2605, -8188, -2178, 6918, 6209, -3305, -8132, -1420, 7308, 5657, -4033, -7992, -586, 7653, 5000, -4774, -7748, 319, 7932, 4231, -5508, -7386, 1284, 8119, 3349, -6211, -6887, 2293, 8190, 2355, -6856, -6240, 3325, 8120, 1259, -7411, -5435, 4352, 7882, 74, -7842, -4469, 5340, 7455, -1177, -8113, -3346, 6250, 6822, -2462, -8189, -2078, 7038, 5971, -3741, -8037, -690, 7656, 4901, -4965, -7628, 782, 8056, 3624, -6077, -6942, 2292, 8190, 2163, -7016, -5972, 3778, 8018, 559, -7718, -4725, 5170, 7509, -1131, -8119, -3227, 6389, 6648, -2834, -8163, -1523, 7352, 5437, -4461, -7808, 318, 7976, 3904, -5913, -7029, 2205, 8190, 2106, -7085, -5827, 4028, 7937, 125, -7873, -4236, 5664, 7186, -1926, -8189, -2325, 6984, 5941, -3912, -7963, -197, 7861, 4243, -5681, -7162, 2007, 8190, 2184, -7075, -5797, 4119, 7894, -105, -7949, -3930, 5957, 6945, -2447, -8182, -1681, 7335, 5371, -4637, -7700, 776, 8089, 3268, -6457, -6491, 3223, 8095, 800, -7699, -4618, 5412, 7295, -1809, -8189, -2227, 7092, 5713, -4289, -7817, 460, 8042, 3467, -6352, -6564, 3157, 8098, 773, -7725, -4514, 5542, 7190, -2074, -8191, -1867, 7293, 5367, -4722, -7629, 1075, 8142, 2807, -6806, -6045, 3934, 7911, -187, -8001, -3595, 6305, 6566, -3215, -8079, -578, 7807, 4234, -5829, -6957, 2583, 8160, 1212, -7599, -4738, 5403, 7238, -2059, -8190, -1716, 7400, 5117, -5052, -7434, 1648, 8187, 2089, -7236, -5385, 4787, 7559, -1360, -8176, -2339, 7120, 5549, -4621, -7629, 1193, 8164, 2463, -7064, -5620, 4556, 7650, -1154, -8164, -2469, 7070, 5596, -4598, -7626, 1238, 8171, 2351, -7140, -5480, 4742, 7552, -1449, -8184, -2113, 7266, 5264, -4987, -7423, 1780, 8190, 1747, -7441, -4943, 5320, 7221, -2233, -8176, -1254, 7642, 4503, -5732, -6934, 2796, 8115, 629, -7852, -3934, 6198, 6534, -3462, -7984, 126, 8036, 3221, -6698, -6004, 4208, 7745, -1006, -8162, -2359, 7191, 5314, -5012, -7368, 1997, 8184, 1340, -7639, -4448, 5833, 6812, -3076, -8057, -176, 7986, 3388, -6626, -6046, 4205, 7727, -1121, -8175, -2134, 7327, 5040, -5332, -7150, 2508, 8138, 695, -7866, -3783, 6384, 6280, -3933, -7814, 890, 8160, 2276, -7279, -5093, 5312, 7141, -2564, -8128, -556, 7914, 3582, -6548, -6080, 4233, 7688, -1317, -8188, -1780, 7516, 4612, -5781, -6785, 3236, 7997, -248, -8090, -2768, 7060, 5389, -5064, -7264, 2379, 8141, 618, -7916, -3524, 6624, 5946, -4454, -7571, 1699, 8188, 1269, -7729, -4064, 6263, 6319, -3992, -7753, 1213, 8187, 1709, -7579, -4406, 6013, 6538, -3700, -7847, 932, 8174, 1940, -7495, -4566, 5898, 6624, -3592, -7874, 858, 8171, 1967, -7493, -4551, 5927, 6585, -3671, -7843, 992, 8180, 1791, -7573, -4359, 6098, 6418, -3935, -7744, 1333, 8190, 1407, -7722, -3983, 6396, 6107, -4372, -7555, 1876, 8173, 812, -7907, -3406, 6793, 5623, -4961, -7238, 2610, 8084, 4, -8084, -2609, 7244, 4934, -5665, -6746, 3512, 7864, -1013, -8186, -1580, 7687, 4003, -6428, -6023, 4539, 7443, -2217, -8135, -314, 8037, 2803, -7172, -5016, 5627, 6744, -3560, -7835, 1167, 8190, 1323, -7790, -3683, 6676, 5696, -4962, -7188, 2807, 8027, -412, -8151, -2012, 7554, 4247, -6301, -6106, 4504, 7427, -2330, -8109, -36, 8098, 2387, -7408, -4530, 6101, 6285, -4296, -7518, 2145, 8130, 169, -8083, -2461, 7386, 4545, -6107, -6263, 4351, 7479, -2264, -8111, 9, 8113, 2234, -7497, -4300, 6315, 6031, -4667, -7305, 2677, 8032, -502, -8169, -1703, 7710, 3772, -6701, -5564, 5217, 6951, -3373, -7845, 1300, 8187, 851, -7965, -2936, 7199, 4809, -5951, -6352, 4308, 7463, -2389, -8077, 321, 8158, 1756, -7713, -3712, 6774, 5420, -5411, -6780, 3713, 7706, -1795, -8153, -227, 8097, 2222, -7551, -4076, 6553, 5675, -5173, -6932, 3493, 7775, -1621, -8166, -337, 8085, 2264, -7548, -4055, 6588, 5609, -5269, -6846, 3666, 7702, -1874, -8138, -11, 8135, 1883, -7703, -3649, 6869, 5213, -5686, -6502, 4217, 7451, -2544, -8022, 751, 8189, 1067, -7954, -2825, 7331, 4434, -6361, -5824, 5093, 6929, -3594, -7706, 1934, 8120, -198, -8164, -1540, 7836, 3196, -7164, -4703, 6178, 5993, -4930, -7018, 3476, 7735, -1886, -8123, 223, 8168, 1436, -7878, -3029, 7267, 4487, -6370, -5759, 5224, 6794, -3882, -7560, 2397, 8029, -831, -8191, -758, 8044, 2306, -7603, -3762, 6884, 5070, -5925, -6190, 4759, 7082, -3436, -7723, 2001, 8093, -509, -8188, -991, 8006, 2447, -7564, -3814, 6876, 5047, -5975, -6113, 4889, 6977, -3660, -7621, 2326, 8026, -932, -8188, -481, 8105, 1868, -7788, -3192, 7246, 4414, -6505, -5505, 5586, 6432, -4522, -7179, 3342, 7726, -2083, -8065, 778, 8190, 536, -8105, -1828, 7814, 3062, -7333, -4213, 6675, 5250, -5863, -6155, 4917, 6906, -3866, -7494, 2733, 7904, -1549, -8137, 340, 8186, 865, -8060, -2044, 7762, 3167, -7307, -4217, 6704, 5169, -5973, -6013, 5128, 6729, -4193, -7310, 3184, 7746, -2127, -8037, 1038, 8176, 57, -8169, -1143, 8017, 2197, -7731, -3205, 7314, 4148, -6783, -5016, 6144, 5793, -5416, -6472, 4609, 7043, -3741, -7503, 2824, 7845, -1877, -8072, 910, 8179, 57, -8174, -1014, 8055, 1946, -7832, -2844, 7507, 3694, -7092, -4489, 6591, 5219, -6017, -5879, 5376, 6460, -4682, -6962, 3941, 7377, -3167, -7709, 2366, 7953, -1551, -8112, 728, 8184, 90, -8176, -898, 8087, 1686, -7925, -2450, 7690, 3180, -7391, -3873, 7030, 4523, -6615, -5127, 6150, 5679, -5644, -6181, 5099, 6626, -4525, -7017, 3923, 7349, -3305, -7626, 2671, 7846, -2031, -8011, 1385, 8121, -743, -8181, 104, 8188, 523, -8149, -1139, 8063, 1736, -7936, -2316, 7768, 2872, -7565, -3405, 7327, 3911, -7060, -4391, 6764, 4840, -6445, -5263, 6104, 5653, -5746, -6015, 5371, 6345, -4986, -6646, 4588, 6916, -4186, -7159, 3776, 7371, -3365, -7558, 2951, 7717, -2540, -7852, 2130, 7960, -1727, -8048, 1327, 8112, -936, -8158, 551, 8182, -178, -8191, -188, 8182, 541, -8160, -884, 8123, 1214, -8075, -1534, 8015, 1839, -7947, -2134, 7868, 2413, -7785, -2682, 7693, 2936, -7599, -3180, 7498, 3408, -7397, -3626, 7292, 3830, -7188, -4024, 7081, 4204, -6978, -4375, 6873, 4532, -6772, -4681, 6672, 4817, -6578, -4945, 6484, 5060, -6398, -5168, 6313, 5265, -6236, -5355, 6163, 5434, -6097, -5506, 6035, 5568, -5981, -5623, 5932, 5669, -5892, -5709, 5857, 5740, -5831, -5765, 5810, 5780, -5798, -5790, 5792, 5791, -5794, -5787, 5803, 5773, -5820, -5754, 5843, 5725, -5874, -5691, 5911, 5647, -5957, -5597, 6007, 5537, -6066, -5471, 6128, 5395, -6199, -5312, 6274, 5217, -6355, -5116, 6440, 5003, -6531, -4883, 6624, 4750, -6722, -4609, 6822, 4455, -6926, -4292, 7029, 4115, -7135, -3929, 7239, 3729, -7345, -3519, 7447, 3295, -7549, -3060, 7646, 2810, -7740, -2550, 7827, 2275, -7909, -1988, 7981, 1688, -8047, -1376, 8100, 1050, -8144, -715, 8173, 365, -8189, -7, 8189, -364, -8173, 742, 8137, -1131, -8083, 1525, 8007, -1928, -7909, 2334, 7787, -2746, -7641, 3157, 7468, -3571, -7269, 3981, 7041, -4388, -6785, 4788, 6499, -5181, -6184, 5560, 5837, -5928, -5462, 6277, 5055, -6608, -4620, 6915, 4154, -7197, -3662, 7449, 3141, -7671, -2597, 7856, 2028, -8005, -1440, 8111, 833, -8175, -212, 8190, -423, -8158, 1063, 8072, -1708, -7936, 2351, 7743, -2990, -7495, 3616, 7189, -4227, -6829, 4815, 6410, -5376, -5937, 5901, 5409, -6389, -4831, 6828, 4203, -7218, -3532, 7548, 2819, -7817, -2072, 8015, 1295, -8142, -496, 8190, -319, -8159, 1139, 8042, -1960, -7842, 2768, 7554, -3558, -7181, 4316, 6721, -5036, -6180, 5704, 5557, -6313, -4863, 6851, 4099, -7311, -3276, 7681, 2400, -7957, -1485, 8128, 537, -8191, 426, 8140, -1395, -7974, 2353, 7688, -3288, -7288, 4181, 6771, -5022, -6146, 5790, 5416, -6476, -4593, 7062, 3685, -7538, -2709, 7890, 1674, -8111, -603, 8190, -491, -8125, 1584, 7910, -2661, -7547, 3695, 7036, -4671, -6388, 5562, 5605, -6354, -4706, 7022, 3702, -7554, -2614, 7932, 1459, -8146, -265, 8183, -946, -8044, 2145, 7721, -3308, -7222, 4403, 6550, -5406, -5721, 6287, 4746, -7026, -3650, 7596, 2453, -7985, -1188, 8173, -120, -8154, 1433, 7921, -2721, -7478, 3944, 6829, -5071, -5991, 6066, 4977, -6900, -3819, 7543, 2540, -7976, -1180, 8176, -226, -8138, 1634, 7853, -3004, -7328, 4290, 6571, -5453, -5604, 6450, 4449, -7249, -3145, 7816, 1727, -8131, -244, 8175, -1260, -7943, 2729, 7435, -4115, -6667, 5364, 5656, -6433, -4438, 7276, 3049, -7860, -1541, 8155, -36, -8149, 1620, 7832, -3154, -7213, 4574, 6308, -5825, -5150, 6852, 3778, -7611, -2246, 8063, 610, -8188, 1058, 7971, -2695, -7417, 4224, 6541, -5584, -5379, 6706, 3972, -7542, -2383, 8045, 675, -8189, 1070, 7959, -2779, -7361, 4367, 6415, -5761, -5161, 6886, 3652, -7689, -1959, 8121, 160, -8157, 1656, 7786, -3401, -7022, 4982, 5896, -6318, -4461, 7333, 2785, -7972, -955, 8190, -937, -7974, 2787, 7324, -4498, -6272, 5968, 4867, -7117, -3184, 7871, 1311, -8185, 645, 8029, -2575, -7409, 4364, 6351, -5907, -4914, 7105, 3174, -7884, -1236, 8187, -789, -7993, 2774, 7300, -4598, -6150, 6140, 4604, -7302, -2758, 8000, 724, -8185, 1365, 7834, -3376, -6967, 5171, 5629, -6631, -3908, 7646, 1911, -8147, 225, 8087, -2357, -7465, 4332, 6314, -6012, -4712, 7270, 2763, -8013, -608, 8175, -1604, -7741, 3705, 6731, -5543, -5216, 6971, 3299, -7881, -1125, 8190, -1147, -7873, 3338, 6939, -5280, -5460, 6813, 3539, -7813, -1330, 8189, -998, -7905, 3252, 6974, -5252, -5466, 6824, 3496, -7836, -1226, 8190, -1159, -7853, 3453, 6841, -5461, -5235, 7003, 3165, -7941, -811, 8180, -1627, -7695, 3928, 6517, -5886, -4746, 7316, 2533, -8084, -81, 8107, -2391, -7378, 4647, 5951, -6476, -3958, 7696, 1578, -8185, 961, 7885, -3419, -6818, 5551, 5077, -7146, -2828, 8037, 288, -8129, 2290, 7399, -4647, -5917, 6538, 3822, -7765, -1326, 8190, -1320, -7764, 3835, 6518, -5956, -4577, 7449, 2139, -8151, 537, 7973, -3167, -6927, 5458, 5116, -7158, -2735, 8069, 38, -8082, 2670, 7184, -5089, -5469, 6934, 3121, -7993, -407, 8130, -2366, -7323, 4870, 5652, -6811, -3310, 7951, 564, -8146, 2257, 7361, -4818, -5684, 6800, 3305, -7958, -514, 8137, -2352, -7308, 4933, 5561, -6906, -3109, 8010, 253, -8101, 2644, 7152, -5212, -5279, 7112, 2712, -8092, 217, 8012, -3128, -6875, 5633, 4817, -7395, -2108, 8167, -895, -7838, 3785, 6438, -6169, -4152, 7709, 1283, -8188, 1771, 7524, -4589, -5804, 6768, 3255, -7996, -238, 8084, -2826, -7013, 5489, 4922, -7366, -2110, 8172, -1022, -7780, 4011, 6234, -6416, -3757, 7868, 707, -8143, 2456, 7185, -5259, -5132, 7265, 2284, -8162, 923, 7797, -3998, -6219, 6456, 3660, -7909, -519, 8114, -2717, -7030, 5526, 4815, -7458, -1820, 8189, -1480, -7592, 4547, 5750, -6879, -2958, 8080, -334, -7944, 3578, 6479, -6234, -3922, 7844, 692, -8130, 2663, 7027, -5573, -4717, 7530, 1583, -8191, 1832, 7423, -4939, -5355, 7184, 2334, -8167, 1107, 7698, -4362, -5853, 6842, 2946, -8095, 499, 7880, -3865, -6228, 6531, 3426, -8003, 15, 7995, -3465, -6499, 6274, 3779, -7914, -342, 8061, -3171, -6679, 6087, 4014, -7847, -572, 8096, -2991, -6779, 5980, 4135, -7811, -676, 8109, -2928, -6807, 5959, 4147, -7812, -653, 8103, -2983, -6764, 6024, 4049, -7851, -504, 8077, -3155, -6647, 6172, 3839, -7920, -228, 8023, -3441, -6448, 6395, 3511, -8010, 175, 7928, -3834, -6156, 6681, 3059, -8101, 703, 7772, -4325, -5756, 7011, 2476, -8171, 1354, 7533, -4897, -5229, 7360, 1754, -8189, 2119, 7183, -5528, -4558, 7694, 893, -8121, 2983, 6693, -6188, -3728, 7975, -106, -7925, 3922, 6031, -6836, -2726, 8154, -1228, -7558, 4900, 5172, -7421, -1552, 8178, -2449, -6979, 5869, 4096, -7883, -217, 7988, -3725, -6149, 6765, 2797, -8152, 1249, 7530, -4997, -5041, 7510, 1288, -8155, 2794, 6752, -6184, -3645, 8016, -395, -7818, 4341, 5621, -7188, -1979, 8190, -2183, -7080, 5787, 4127, -7895, -93, 7941, -3976, -5902, 7005, 2298, -8189, 1921, 7196, -5639, -4280, 7854, 207, -7962, 3929, 5916, -7011, -2261, 8190, -2021, -7132, 5756, 4111, -7916, 49, 7888, -4207, -5669, 7200, 1860, -8185, 2477, 6869, -6127, -3612, 8048, -680, -7686, 4784, 5125, -7529, -1089, 8112, -3271, -6353, 6690, 2745, -8172, 1670, 7267, -5607, -4228, 7900, -66, -7864, 4347, 5492, -7346, -1479, 8153, -2987, -6516, 6562, 2909, -8162, 1585, 7287, -5607, -4189, 7923, -199, -7813, 4533, 5293, -7477, -1131, 8106, -3393, -6211, 6864, 2367, -8191, 2227, 6938, -6129, -3490, 8093, -1076, -7486, 5306, 4482, -7845, -34, 7863, -4435, -5341, 7474, 1078, -8090, 3542, 6062, -7014, -2044, 8184, -2658, -6657, 6487, 2917, -8171, 1798, 7129, -5924, -3699, 8066, -984, -7495, 5341, 4384, -7897, 222, 7765, -4762, -4979, 7677, 476, -7957, 4198, 5486, -7429, -1108, 8081, -3666, -5914, 7164, 1668, -8154, 3171, 6267, -6900, -2160, 8185, -2725, -6558, 6644, 2580, -8190, 2330, 6790, -6411, -2934, 8176, -1994, -6973, 6203, 3221, -8153, 1716, 7111, -6032, -3447, 8126, -1501, -7213, 5898, 3610, -8105, 1346, 7278, -5808, -3716, 8088, -1257, -7315, 5761, 3761, -8083, 1230, 7320, -5761, -3751, 8086, -1269, -7298, 5806, 3681, -8100, 1370, 7243, -5897, -3555, 8121, -1536, -7158, 6029, 3367, -8148, 1762, 7035, -6201, -3119, 8171, -2052, -6872, 6406, 2806, -8189, 2399, 6660, -6641, -2427, 8188, -2804, -6396, 6895, 1978, -8164, 3259) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L21_i
    );

    L21C31_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-5500, -7516, 672, 7947, 4422, -5116, -7697, 195, 7822, 4796, -4766, -7833, -218, 7694, 5104, -4457, -7931, -566, 7573, 5353, -4194, -8000, -849, 7465, 5545, -3981, -8047, -1067, 7378, 5686, -3823, -8076, -1220, 7316, 5778, -3720, -8093, -1309, 7281, 5823, -3674, -8099, -1334, 7275, 5823, -3686, -8095, -1295, 7299, 5777, -3756, -8080, -1192, 7351, 5684, -3882, -8053, -1025, 7429, 5543, -4063, -8010, -793, 7530, 5349, -4297, -7946, -496, 7646, 5100, -4580, -7853, -134, 7773, 4790, -4908, -7726, 293, 7900, 4416, -5273, -7553, 784, 8018, 3971, -5667, -7326, 1335, 8115, 3452, -6082, -7034, 1944, 8177, 2855, -6504, -6666, 2603, 8188, 2178, -6918, -6211, 3302, 8131, 1421, -7308, -5659, 4031, 7991, 587, -7654, -5002, 4772, 7748, -318, -7932, -4233, 5506, 7385, -1283, -8120, -3351, 6209, 6887, -2293, -8191, -2358, 6854, 6240, -3325, -8121, -1261, 7409, 5435, -4352, -7883, -76, 7840, 4469, -5340, -7457, 1175, 8112, 3346, -6250, -6823, 2459, 8188, 2079, -7039, -5973, 3738, 8036, 691, -7657, -4904, 4962, 7627, -782, -8057, -3626, 6075, 6942, -2291, -8191, -2166, 7014, 5972, -3778, -8020, -561, 7716, 4726, -5170, -7511, 1129, 8118, 3227, -6389, -6649, 2832, 8162, 1523, -7352, -5439, 4459, 7807, -317, -7977, -3907, 5911, 7028, -2204, -8191, -2108, 7083, 5827, -4028, -7939, -127, 7872, 4237, -5664, -7188, 1924, 8188, 2325, -6984, -5943, 3910, 7962, 198, -7862, -4246, 5679, 7162, -2006, -8191, -2186, 7074, 5797, -4119, -7896, 102, 7948, 3930, -5957, -6947, 2444, 8181, 1681, -7335, -5373, 4635, 7700, -776, -8089, -3271, 6455, 6491, -3222, -8096, -802, 7697, 4619, -5412, -7296, 1807, 8188, 2227, -7093, -5715, 4287, 7816, -460, -8043, -3470, 6350, 6563, -3157, -8099, -775, 7723, 4514, -5542, -7192, 2072, 8190, 1868, -7294, -5369, 4720, 7628, -1074, -8143, -2809, 6805, 6045, -3934, -7913, 185, 8000, 3595, -6305, -6568, 3213, 8078, 579, -7808, -4236, 5827, 6957, -2583, -8161, -1214, 7597, 4738, -5403, -7240, 2057, 8189, 1716, -7400, -5119, 5050, 7433, -1648, -8188, -2091, 7235, 5385, -4787, -7560, 1358, 8175, 2339, -7120, -5551, 4619, 7629, -1193, -8165, -2465, 7062, 5620, -4556, -7651, 1152, 8163, 2469, -7070, -5598, 4596, 7626, -1238, -8171, -2353, 7139, 5480, -4742, -7553, 1446, 8183, 2113, -7267, -5266, 4985, 7422, -1780, -8191, -1749, 7439, 4943, -5320, -7223, 2231, 8175, 1254, -7643, -4505, 5730, 6933, -2796, -8116, -631, 7850, 3934, -6199, -6536, 3460, 7983, -125, -8037, -3223, 6696, 6003, -4208, -7747, 1004, 8161, 2359, -7191, -5316, 5010, 7368, -1997, -8185, -1343, 7638, 4448, -5833, -6814, 3074, 8056, 176, -7987, -3390, 6625, 6046, -4205, -7728, 1119, 8174, 2134, -7327, -5042, 5330, 7149, -2508, -8139, -697, 7865, 3783, -6384, -6281, 3931, 7814, -890, -8161, -2278, 7278, 5093, -5312, -7142, 2562, 8127, 556, -7915, -3584, 6546, 6079, -4233, -7689, 1315, 8187, 1780, -7516, -4614, 5780, 6785, -3236, -7998, 245, 8089, 2768, -7061, -5391, 5062, 7264, -2379, -8143, -620, 7914, 3524, -6625, -5948, 4453, 7570, -1699, -8189, -1271, 7728, 4064, -6263, -6321, 3990, 7752, -1213, -8188, -1711, 7577, 4406, -6014, -6540, 3698, 7846, -932, -8175, -1942, 7494, 4566, -5899, -6626, 3590, 7873, -858, -8172, -1969, 7492, 4550, -5928, -6587, 3669, 7842, -992, -8181, -1793, 7572, 4359, -6098, -6420, 3933, 7743, -1333, -8191, -1409, 7720, 3983, -6396, -6108, 4370, 7554, -1876, -8174, -814, 7906, 3405, -6793, -5625, 4959, 7238, -2610, -8085, -6, 8082, 2609, -7245, -4935, 5663, 6745, -3512, -7865, 1011, 8185, 1579, -7688, -4005, 6427, 6023, -4540, -7444, 2215, 8134, 314, -8038, -2804, 7170, 5016, -5627, -6746, 3558, 7834, -1167, -8191, -1325, 7789, 3683, -6676, -5698, 4961, 7188, -2807, -8029, 410, 8150, 2012, -7555, -4249, 6299, 6105, -4504, -7428, 2328, 8108, 36, -8099, -2388, 7407, 4529, -6101, -6287, 4295, 7517, -2146, -8131, -171, 8082, 2461, -7387, -4547, 6106, 6262, -4351, -7480, 2262, 8110, -9, -8114, -2236, 7496, 4300, -6316, -6032, 4666, 7305, -2678, -8033, 500, 8168, 1702, -7711, -3774, 6699, 5564, -5217, -6952, 3372, 7845, -1301, -8188, -853, 7964, 2936, -7199, -4811, 5949, 6352, -4308, -7464, 2388, 8076, -321, -8159, -1758, 7712, 3712, -6775, -5422, 5410, 6779, -3714, -7707, 1793, 8152, 226, -8098, -2224, 7550, 4076, -6554, -5676, 5171, 6931, -3494, -7777, 1619, 8165, 337, -8086, -2266, 7546, 4055, -6588, -5610, 5268, 6846, -3666, -7703, 1872, 8137, 11, -8136, -1885, 7702, 3648, -6870, -5214, 5685, 6501, -4217, -7452, 2543, 8021, -752, -8190, -1068, 7953, 2824, -7332, -4435, 6360, 5823, -5093, -6930, 3592, 7705, -1935, -8121, 196, 8163, 1539, -7837, -3197, 7163, 4702, -6178, -5994, 4929, 7017, -3477, -7736, 1884, 8122, -224, -8169, -1438, 7877, 3028, -7268, -4489, 6369, 5759, -5224, -6795, 3881, 7559, -2397, -8030, 830, 8190, 757, -8045, -2308, 7601, 3762, -6885, -5072, 5924, 6189, -4760, -7083, 3435, 7723, -2002, -8094, 508, 8187, 991, -8007, -2448, 7563, 3814, -6877, -5049, 5974, 6112, -4890, -6978, 3659, 7620, -2326, -8027, 931, 8187, 480, -8106, -1869, 7786, 3192, -7247, -4416, 6504, 5504, -5587, -6434, 4521, 7178, -3343, -7727, 2082, 8064, -778, -8191, -538, 8104, 1827, -7815, -3063, 7332, 4212, -6676, -5251, 5862, 6154, -4918, -6908, 3864, 7493, -2733, -7906, 1548, 8136, -340, -8187, -867, 8059, 2043, -7763, -3168, 7306, 4216, -6705, -5171, 5971, 6012, -5128, -6730, 4191, 7309, -3185, -7748, 2125, 8036, -1039, -8177, -58, 8168, 1142, -8018, -2198, 7730, 3205, -7315, -4150, 6782, 5015, -6145, -5794, 5415, 6471, -4609, -7044, 3739, 7502, -2824, -7846, 1875, 8071, -911, -8180, -58, 8173, 1014, -8056, -1948, 7831, 2844, -7508, -3695, 7091, 4489, -6592, -5220, 6016, 5878, -5377, -6461, 4681, 6961, -3942, -7379, 3166, 7708, -2366, -7954, 1550, 8111, -729, -8185, -91, 8175, 898, -8088, -1687, 7924, 2449, -7691, -3181, 7390, 3873, -7030, -4524, 6614, 5126, -6151, -5680, 5643, 6180, -5099, -6627, 4523, 7016, -3924, -7350, 3304, 7626, -2672, -7847, 2030, 8010, -1386, -8122, 741, 8180, -105, -8189, -524, 8148, 1138, -8064, -1737, 7935, 2315, -7769, -2873, 7564, 3404, -7328, -3912, 7059, 4390, -6765, -4842, 6444, 5262, -6105, -5654, 5745, 6014, -5372, -6346, 4985, 6645, -4589, -6917, 4184, 7158, -3776, -7372, 3364, 7557, -2952, -7718, 2539, 7851, -2131, -7961, 1726, 8047, -1328, -8113, 935, 8157, -552, -8183, 177, 8190, 187, -8183, -542, 8159, 884, -8124, -1215, 8074, 1533, -8016, -1840, 7946, 2133, -7869, -2414, 7784, 2681, -7694, -2937, 7598, 3179, -7499, -3409, 7396, 3626, -7293, -3831, 7187, 4023, -7082, -4205, 6976, 4374, -6874, -4534, 6771, 4680, -6673, -4818, 6577, 4944, -6485, -5061, 6397, 5167, -6314, -5266, 6235, 5354, -6164, -5435, 6096, 5505, -6036, -5569, 5980, 5622, -5933, -5670, 5891, 5708, -5858, -5741, 5830, 5764, -5811, -5781, 5797, 5789, -5793, -5792, 5793, 5786, -5804, -5774, 5819, 5753, -5844, -5726, 5873, 5690, -5912, -5648, 5956, 5596, -6008, -5538, 6065, 5470, -6129, -5396, 6198, 5311, -6275, -5218, 6354, 5115, -6441, -5004, 6530, 4882, -6625, -4751, 6722, 4608, -6823, -4456, 6925, 4291, -7030, -4116, 7134, 3928, -7240, -3730, 7344, 3518, -7449, -3296, 7548, 3059, -7647, -2811, 7739, 2549, -7828, -2276, 7908, 1987, -7982, -1689, 8046, 1375, -8101, -1051, 8143, 713, -8174, -366, 8188, 6, -8190, 363, 8172, -743, -8138, 1130, 8082, -1527, -8008, 1927, 7908, -2335, -7788, 2745, 7640, -3158, -7469, 3570, 7268, -3982, -7042, 4387, 6784, -4789, -6500, 5180, 6183, -5561, -5838, 5927, 5461, -6278, -5056, 6607, 4619, -6916, -4155, 7197, 3661, -7451, -3142, 7671, 2596, -7858, -2029, 8004, 1439, -8112, -833, 8174, 210, -8191, 422, 8157, -1064, -8073, 1708, 7935, -2352, -7743, 2989, 7494, -3617, -7190, 4226, 6828, -4816, -6411, 5375, 5936, -5903, -5410, 6388, 4830, -6830, -4204, 7217, 3531, -7549, -2819, 7816, 2071, -8016, -1295, 8141, 495, -8191, 318, 8158, -1140, -8043, 1959, 7841, -2769, -7555, 3558, 7180, -4318, -6721, 5035, 6178, -5705, -5558, 6313, 4862, -6852, -4099, 7310, 3275, -7682, -2401, 7956, 1483, -8129, -538, 8190, -427, -8141, 1394, 7973, -2354, -7689, 3287, 7287, -4182, -6772, 5021, 6145, -5791, -5416, 6476, 4592, -7063, -3686, 7538, 2707, -7891, -1675, 8110, 602, -8191, 490, 8124, -1586, -7911, 2660, 7546, -3697, -7037, 4670, 6386, -5564, -5606, 6353, 4705, -7023, -3702, 7554, 2612, -7933, -1460, 8145, 264, -8184, 946, 8043, -2147, -7722, 3307, 7221, -4404, -6551, 5405, 5720, -6288, -4747, 7025, 3649, -7598, -2454, 7984, 1186, -8174, 120, 8153, -1435, -7922, 2720, 7477, -3945, -6830, 5071, 5989, -6067, -4978, 6899, 3817, -7544, -2541, 7975, 1179, -8177, 225, 8137, -1635, -7854, 3003, 7327, -4291, -6572, 5453, 5602, -6452, -4450, 7249, 3144, -7817, -1728, 8130, 242, -8176, 1259, 7942, -2730, -7436, 4115, 6665, -5366, -5656, 6433, 4436, -7277, -3050, 7859, 1540, -8156, 36, 8148, -1621, -7833, 3153, 7212, -4575, -6309, 5825, 5149, -6853, -3778, 7610, 2244, -8065, -611, 8187, -1060, -7972, 2694, 7416, -4226, -6542, 5583, 5377, -6708, -3972, 7541, 2381, -8046, -676, 8188, -1072, -7960, 2779, 7360, -4369, -6415, 5760, 5160, -6888, -3652, 7688, 1958, -8122, -160, 8156, -1658, -7786, 3401, 7021, -4983, -5896, 6318, 4460, -7334, -2786, 7971, 954, -8191, 937, 7973, -2789, -7325, 4497, 6271, -5970, -4867, 7117, 3182, -7872, -1311, 8184, -646, -8030, 2575, 7408, -4365, -6351, 5906, 4912, -7106, -3174, 7883, 1234, -8188, 789, 7991, -2776, -7301, 4598, 6148, -6142, -4604, 7301, 2757, -8001, -725, 8184, -1366, -7835, 3376, 6965, -5173, -5629, 6630, 3906, -7648, -1911, 8146, -226, -8087, 2356, 7464, -4333, -6315, 6012, 4710, -7271, -2764, 8012, 606, -8176, 1603, 7740, -3707, -6732, 5542, 5214, -6973, -3300, 7880, 1123, -8191, 1147, 7871, -3340, -6940, 5280, 5458, -6815, -3540, 7812, 1328, -8190, 997, 7904, -3254, -6974, 5252, 5464, -6826, -3496, 7835, 1224, -8191, 1158, 7852, -3454, -6841, 5461, 5234, -7004, -3166, 7940, 809, -8181, 1627, 7694, -3929, -6517, 5885, 4744, -7317, -2533, 8083, 79, -8108, 2391, 7376, -4649, -5952, 6476, 3957, -7697, -1578, 8185, -963, -7886, 3419, 6817, -5553, -5077, 7146, 2827, -8038, -288, 8128, -2291, -7400, 4647, 5916, -6539, -3822, 7764, 1324, -8191, 1320, 7763, -3836, -6518, 5956, 4576, -7451, -2139, 8150, -539, -7973, 3167, 6926, -5460, -5117, 7158, 2733, -8070, -39, 8081, -2672, -7184, 5088, 5467, -6936, -3121, 7992, 405, -8131, 2365, 7322, -4871, -5653, 6811, 3308, -7952, -564, 8145, -2259, -7362, 4818, 5682, -6802, -3305, 7957, 512, -8138, 2352, 7307, -4935, -5561, 6905, 3107, -8011, -253, 8100, -2646, -7153, 5211, 5277, -7113, -2712, 8092, -218, -8013, 3128, 6873, -5634, -4817, 7395, 2106, -8168, 895, 7837, -3787, -6438, 6168, 4150, -7710, -1283, 8187, -1773, -7525, 4589, 5802, -6770, -3255, 7995, 236, -8085, 2826, 7011, -5491, -4922, 7366, 2108, -8173, 1022, 7779, -4013, -6235, 6416, 3755, -7869, -707, 8142, -2458, -7185, 5259, 5130, -7266, -2284, 8161, -925, -7798, 3998, 6217, -6458, -3660, 7908, 517, -8114, 2717, 7028, -5528, -4815, 7457, 1818, -8190, 1480, 7591, -4549, -5750, 6879, 2956, -8081, 334, 7943, -3580, -6479, 6233, 3920, -7845, -692, 8128, -2665, -7027, 5573, 4715, -7532, -1583, 8190, -1834, -7424, 4939, 5353, -7186, -2334, 8166, -1109, -7699, 4362, 5851, -6843, -2946, 8094, -501, -7881, 3865, 6226, -6533, -3426, 8002, -17, -7995, 3465, 6497, -6276, -3779, 7914, 340, -8062, 3171, 6677, -6089, -4014, 7846, 570, -8097, 2991, 6778, -5982, -4135, 7810, 674, -8110, 2928, 6805, -5961, -4147, 7812, 651, -8104, 2983, 6762, -6026, -4049, 7850, 502, -8078, 3155, 6645, -6174, -3839, 7920, 226, -8024, 3441, 6447, -6397, -3511, 8009, -177, -7928, 3834, 6155, -6683, -3059, 8100, -706, -7773, 4325, 5754, -7013, -2475, 8170, -1357, -7534, 4897, 5227, -7361, -1754, 8188, -2122, -7184, 5528, 4556, -7696, -892, 8119, -2985, -6693, 6188, 3726, -7976, 106, 7923, -3924, -6031, 6835, 2724, -8155, 1228, 7557, -4902, -5172, 7421, 1550, -8178, 2449, 6977, -5871, -4096, 7882, 215, -7989, 3725, 6147, -6766, -2797, 8151, -1251, -7530, 4997, 5039, -7511, -1288, 8153, -2796, -6752, 6184, 3643, -8018, 395, 7816, -4343, -5621, 7187, 1977, -8191, 2184, 7078, -5789, -4127, 7894, 91, -7941, 3976, 5900, -7007, -2298, 8188, -1923, -7196, 5639, 4278, -7855, -207, 7961, -3931, -5916, 7011, 2258, -8191, 2022, 7131, -5758, -4111, 7915, -52, -7889, 4208, 5667, -7202, -1860, 8184, -2479, -6869, 6127, 3609, -8049, 680, 7684, -4787, -5125, 7529, 1087, -8113, 3271, 6351, -6692, -2744, 8171, -1672, -7267, 5607, 4226, -7901, 66, 7863, -4350, -5492, 7346, 1477, -8154, 2987, 6514, -6564, -2908, 8162, -1587, -7287, 5607, 4187, -7924, 199, 7811, -4535, -5293, 7477, 1128, -8106, 3393, 6209, -6866, -2366, 8190, -2229, -6939, 6129, 3488, -8094, 1077, 7484, -5308, -4482, 7845, 32, -7863, 4435, 5338, -7476, -1078, 8089, -3545, -6062, 7014, 2041, -8185, 2658, 6655, -6489, -2917, 8170, -1801, -7129, 5924, 3697, -8068, 984, 7494, -5343, -4384, 7896, -224, -7766, 4763, 4977, -7679, -475, 7956, -4201, -5485, 7429, 1105, -8081, 3666, 5912, -7166, -1667, 8153, -3174, -6267, 6900, 2157, -8186, 2726, 6556, -6646, -2579, 8189, -2333, -6790, 6411, 2932, -8177, 1995, 6971, -6205, -3221, 8152, -1718, -7111, 6032, 3445, -8128, 1501, 7211, -5900, -3610, 8104, -1349, -7278, 5808, 3713, -8089, 1258, 7313, -5763, -3761, 8082, -1233, -7320, 5762, 3749, -8087, 1270, 7296, -5808, -3681, 8100, -1372, -7243, 5897, 3553, -8122, 1536, 7156, -6031, -3367, 8147, -1765, -7035, 6201, 3117, -8172, 2052, 6870, -6408, -2805, 8188, -2401, -6660, 6641, 2425, -8189, 2804, 6394, -6897, -1978, 8163, -3261) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L21C31_i
    );

    L21C32_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (5500, 7514, -675, -7949, -4422, 5117, 7696, -198, -7824, -4795, 4767, 7831, 215, -7696, -5104, 4457, 7929, 564, -7574, -5352, 4194, 7999, 846, -7467, -5545, 3982, 8045, 1064, -7380, -5686, 3823, 8075, 1217, -7317, -5778, 3720, 8092, 1306, -7282, -5823, 3675, 8098, 1331, -7277, -5823, 3687, 8093, 1292, -7300, -5777, 3756, 8079, 1190, -7353, -5684, 3883, 8052, 1023, -7431, -5542, 4064, 8009, 791, -7531, -5349, 4298, 7944, 494, -7648, -5100, 4581, 7852, 132, -7774, -4790, 4908, 7724, -296, -7902, -4415, 5273, 7552, -786, -8020, -3971, 5667, 7325, -1338, -8116, -3452, 6082, 7032, -1946, -8178, -2855, 6504, 6664, -2605, -8188, -2178, 6918, 6209, -3305, -8132, -1420, 7308, 5657, -4033, -7992, -586, 7653, 5000, -4774, -7748, 319, 7932, 4231, -5508, -7386, 1284, 8119, 3349, -6211, -6887, 2293, 8190, 2355, -6856, -6240, 3325, 8120, 1259, -7411, -5435, 4352, 7882, 74, -7842, -4469, 5340, 7455, -1177, -8113, -3346, 6250, 6822, -2462, -8189, -2078, 7038, 5971, -3741, -8037, -690, 7656, 4901, -4965, -7628, 782, 8056, 3624, -6077, -6942, 2292, 8190, 2163, -7016, -5972, 3778, 8018, 559, -7718, -4725, 5170, 7509, -1131, -8119, -3227, 6389, 6648, -2834, -8163, -1523, 7352, 5437, -4461, -7808, 318, 7976, 3904, -5913, -7029, 2205, 8190, 2106, -7085, -5827, 4028, 7937, 125, -7873, -4236, 5664, 7186, -1926, -8189, -2325, 6984, 5941, -3912, -7963, -197, 7861, 4243, -5681, -7162, 2007, 8190, 2184, -7075, -5797, 4119, 7894, -105, -7949, -3930, 5957, 6945, -2447, -8182, -1681, 7335, 5371, -4637, -7700, 776, 8089, 3268, -6457, -6491, 3223, 8095, 800, -7699, -4618, 5412, 7295, -1809, -8189, -2227, 7092, 5713, -4289, -7817, 460, 8042, 3467, -6352, -6564, 3157, 8098, 773, -7725, -4514, 5542, 7190, -2074, -8191, -1867, 7293, 5367, -4722, -7629, 1075, 8142, 2807, -6806, -6045, 3934, 7911, -187, -8001, -3595, 6305, 6566, -3215, -8079, -578, 7807, 4234, -5829, -6957, 2583, 8160, 1212, -7599, -4738, 5403, 7238, -2059, -8190, -1716, 7400, 5117, -5052, -7434, 1648, 8187, 2089, -7236, -5385, 4787, 7559, -1360, -8176, -2339, 7120, 5549, -4621, -7629, 1193, 8164, 2463, -7064, -5620, 4556, 7650, -1154, -8164, -2469, 7070, 5596, -4598, -7626, 1238, 8171, 2351, -7140, -5480, 4742, 7552, -1449, -8184, -2113, 7266, 5264, -4987, -7423, 1780, 8190, 1747, -7441, -4943, 5320, 7221, -2233, -8176, -1254, 7642, 4503, -5732, -6934, 2796, 8115, 629, -7852, -3934, 6198, 6534, -3462, -7984, 126, 8036, 3221, -6698, -6004, 4208, 7745, -1006, -8162, -2359, 7191, 5314, -5012, -7368, 1997, 8184, 1340, -7639, -4448, 5833, 6812, -3076, -8057, -176, 7986, 3388, -6626, -6046, 4205, 7727, -1121, -8175, -2134, 7327, 5040, -5332, -7150, 2508, 8138, 695, -7866, -3783, 6384, 6280, -3933, -7814, 890, 8160, 2276, -7279, -5093, 5312, 7141, -2564, -8128, -556, 7914, 3582, -6548, -6080, 4233, 7688, -1317, -8188, -1780, 7516, 4612, -5781, -6785, 3236, 7997, -248, -8090, -2768, 7060, 5389, -5064, -7264, 2379, 8141, 618, -7916, -3524, 6624, 5946, -4454, -7571, 1699, 8188, 1269, -7729, -4064, 6263, 6319, -3992, -7753, 1213, 8187, 1709, -7579, -4406, 6013, 6538, -3700, -7847, 932, 8174, 1940, -7495, -4566, 5898, 6624, -3592, -7874, 858, 8171, 1967, -7493, -4551, 5927, 6585, -3671, -7843, 992, 8180, 1791, -7573, -4359, 6098, 6418, -3935, -7744, 1333, 8190, 1407, -7722, -3983, 6396, 6107, -4372, -7555, 1876, 8173, 812, -7907, -3406, 6793, 5623, -4961, -7238, 2610, 8084, 4, -8084, -2609, 7244, 4934, -5665, -6746, 3512, 7864, -1013, -8186, -1580, 7687, 4003, -6428, -6023, 4539, 7443, -2217, -8135, -314, 8037, 2803, -7172, -5016, 5627, 6744, -3560, -7835, 1167, 8190, 1323, -7790, -3683, 6676, 5696, -4962, -7188, 2807, 8027, -412, -8151, -2012, 7554, 4247, -6301, -6106, 4504, 7427, -2330, -8109, -36, 8098, 2387, -7408, -4530, 6101, 6285, -4296, -7518, 2145, 8130, 169, -8083, -2461, 7386, 4545, -6107, -6263, 4351, 7479, -2264, -8111, 9, 8113, 2234, -7497, -4300, 6315, 6031, -4667, -7305, 2677, 8032, -502, -8169, -1703, 7710, 3772, -6701, -5564, 5217, 6951, -3373, -7845, 1300, 8187, 851, -7965, -2936, 7199, 4809, -5951, -6352, 4308, 7463, -2389, -8077, 321, 8158, 1756, -7713, -3712, 6774, 5420, -5411, -6780, 3713, 7706, -1795, -8153, -227, 8097, 2222, -7551, -4076, 6553, 5675, -5173, -6932, 3493, 7775, -1621, -8166, -337, 8085, 2264, -7548, -4055, 6588, 5609, -5269, -6846, 3666, 7702, -1874, -8138, -11, 8135, 1883, -7703, -3649, 6869, 5213, -5686, -6502, 4217, 7451, -2544, -8022, 751, 8189, 1067, -7954, -2825, 7331, 4434, -6361, -5824, 5093, 6929, -3594, -7706, 1934, 8120, -198, -8164, -1540, 7836, 3196, -7164, -4703, 6178, 5993, -4930, -7018, 3476, 7735, -1886, -8123, 223, 8168, 1436, -7878, -3029, 7267, 4487, -6370, -5759, 5224, 6794, -3882, -7560, 2397, 8029, -831, -8191, -758, 8044, 2306, -7603, -3762, 6884, 5070, -5925, -6190, 4759, 7082, -3436, -7723, 2001, 8093, -509, -8188, -991, 8006, 2447, -7564, -3814, 6876, 5047, -5975, -6113, 4889, 6977, -3660, -7621, 2326, 8026, -932, -8188, -481, 8105, 1868, -7788, -3192, 7246, 4414, -6505, -5505, 5586, 6432, -4522, -7179, 3342, 7726, -2083, -8065, 778, 8190, 536, -8105, -1828, 7814, 3062, -7333, -4213, 6675, 5250, -5863, -6155, 4917, 6906, -3866, -7494, 2733, 7904, -1549, -8137, 340, 8186, 865, -8060, -2044, 7762, 3167, -7307, -4217, 6704, 5169, -5973, -6013, 5128, 6729, -4193, -7310, 3184, 7746, -2127, -8037, 1038, 8176, 57, -8169, -1143, 8017, 2197, -7731, -3205, 7314, 4148, -6783, -5016, 6144, 5793, -5416, -6472, 4609, 7043, -3741, -7503, 2824, 7845, -1877, -8072, 910, 8179, 57, -8174, -1014, 8055, 1946, -7832, -2844, 7507, 3694, -7092, -4489, 6591, 5219, -6017, -5879, 5376, 6460, -4682, -6962, 3941, 7377, -3167, -7709, 2366, 7953, -1551, -8112, 728, 8184, 90, -8176, -898, 8087, 1686, -7925, -2450, 7690, 3180, -7391, -3873, 7030, 4523, -6615, -5127, 6150, 5679, -5644, -6181, 5099, 6626, -4525, -7017, 3923, 7349, -3305, -7626, 2671, 7846, -2031, -8011, 1385, 8121, -743, -8181, 104, 8188, 523, -8149, -1139, 8063, 1736, -7936, -2316, 7768, 2872, -7565, -3405, 7327, 3911, -7060, -4391, 6764, 4840, -6445, -5263, 6104, 5653, -5746, -6015, 5371, 6345, -4986, -6646, 4588, 6916, -4186, -7159, 3776, 7371, -3365, -7558, 2951, 7717, -2540, -7852, 2130, 7960, -1727, -8048, 1327, 8112, -936, -8158, 551, 8182, -178, -8191, -188, 8182, 541, -8160, -884, 8123, 1214, -8075, -1534, 8015, 1839, -7947, -2134, 7868, 2413, -7785, -2682, 7693, 2936, -7599, -3180, 7498, 3408, -7397, -3626, 7292, 3830, -7188, -4024, 7081, 4204, -6978, -4375, 6873, 4532, -6772, -4681, 6672, 4817, -6578, -4945, 6484, 5060, -6398, -5168, 6313, 5265, -6236, -5355, 6163, 5434, -6097, -5506, 6035, 5568, -5981, -5623, 5932, 5669, -5892, -5709, 5857, 5740, -5831, -5765, 5810, 5780, -5798, -5790, 5792, 5791, -5794, -5787, 5803, 5773, -5820, -5754, 5843, 5725, -5874, -5691, 5911, 5647, -5957, -5597, 6007, 5537, -6066, -5471, 6128, 5395, -6199, -5312, 6274, 5217, -6355, -5116, 6440, 5003, -6531, -4883, 6624, 4750, -6722, -4609, 6822, 4455, -6926, -4292, 7029, 4115, -7135, -3929, 7239, 3729, -7345, -3519, 7447, 3295, -7549, -3060, 7646, 2810, -7740, -2550, 7827, 2275, -7909, -1988, 7981, 1688, -8047, -1376, 8100, 1050, -8144, -715, 8173, 365, -8189, -7, 8189, -364, -8173, 742, 8137, -1131, -8083, 1525, 8007, -1928, -7909, 2334, 7787, -2746, -7641, 3157, 7468, -3571, -7269, 3981, 7041, -4388, -6785, 4788, 6499, -5181, -6184, 5560, 5837, -5928, -5462, 6277, 5055, -6608, -4620, 6915, 4154, -7197, -3662, 7449, 3141, -7671, -2597, 7856, 2028, -8005, -1440, 8111, 833, -8175, -212, 8190, -423, -8158, 1063, 8072, -1708, -7936, 2351, 7743, -2990, -7495, 3616, 7189, -4227, -6829, 4815, 6410, -5376, -5937, 5901, 5409, -6389, -4831, 6828, 4203, -7218, -3532, 7548, 2819, -7817, -2072, 8015, 1295, -8142, -496, 8190, -319, -8159, 1139, 8042, -1960, -7842, 2768, 7554, -3558, -7181, 4316, 6721, -5036, -6180, 5704, 5557, -6313, -4863, 6851, 4099, -7311, -3276, 7681, 2400, -7957, -1485, 8128, 537, -8191, 426, 8140, -1395, -7974, 2353, 7688, -3288, -7288, 4181, 6771, -5022, -6146, 5790, 5416, -6476, -4593, 7062, 3685, -7538, -2709, 7890, 1674, -8111, -603, 8190, -491, -8125, 1584, 7910, -2661, -7547, 3695, 7036, -4671, -6388, 5562, 5605, -6354, -4706, 7022, 3702, -7554, -2614, 7932, 1459, -8146, -265, 8183, -946, -8044, 2145, 7721, -3308, -7222, 4403, 6550, -5406, -5721, 6287, 4746, -7026, -3650, 7596, 2453, -7985, -1188, 8173, -120, -8154, 1433, 7921, -2721, -7478, 3944, 6829, -5071, -5991, 6066, 4977, -6900, -3819, 7543, 2540, -7976, -1180, 8176, -226, -8138, 1634, 7853, -3004, -7328, 4290, 6571, -5453, -5604, 6450, 4449, -7249, -3145, 7816, 1727, -8131, -244, 8175, -1260, -7943, 2729, 7435, -4115, -6667, 5364, 5656, -6433, -4438, 7276, 3049, -7860, -1541, 8155, -36, -8149, 1620, 7832, -3154, -7213, 4574, 6308, -5825, -5150, 6852, 3778, -7611, -2246, 8063, 610, -8188, 1058, 7971, -2695, -7417, 4224, 6541, -5584, -5379, 6706, 3972, -7542, -2383, 8045, 675, -8189, 1070, 7959, -2779, -7361, 4367, 6415, -5761, -5161, 6886, 3652, -7689, -1959, 8121, 160, -8157, 1656, 7786, -3401, -7022, 4982, 5896, -6318, -4461, 7333, 2785, -7972, -955, 8190, -937, -7974, 2787, 7324, -4498, -6272, 5968, 4867, -7117, -3184, 7871, 1311, -8185, 645, 8029, -2575, -7409, 4364, 6351, -5907, -4914, 7105, 3174, -7884, -1236, 8187, -789, -7993, 2774, 7300, -4598, -6150, 6140, 4604, -7302, -2758, 8000, 724, -8185, 1365, 7834, -3376, -6967, 5171, 5629, -6631, -3908, 7646, 1911, -8147, 225, 8087, -2357, -7465, 4332, 6314, -6012, -4712, 7270, 2763, -8013, -608, 8175, -1604, -7741, 3705, 6731, -5543, -5216, 6971, 3299, -7881, -1125, 8190, -1147, -7873, 3338, 6939, -5280, -5460, 6813, 3539, -7813, -1330, 8189, -998, -7905, 3252, 6974, -5252, -5466, 6824, 3496, -7836, -1226, 8190, -1159, -7853, 3453, 6841, -5461, -5235, 7003, 3165, -7941, -811, 8180, -1627, -7695, 3928, 6517, -5886, -4746, 7316, 2533, -8084, -81, 8107, -2391, -7378, 4647, 5951, -6476, -3958, 7696, 1578, -8185, 961, 7885, -3419, -6818, 5551, 5077, -7146, -2828, 8037, 288, -8129, 2290, 7399, -4647, -5917, 6538, 3822, -7765, -1326, 8190, -1320, -7764, 3835, 6518, -5956, -4577, 7449, 2139, -8151, 537, 7973, -3167, -6927, 5458, 5116, -7158, -2735, 8069, 38, -8082, 2670, 7184, -5089, -5469, 6934, 3121, -7993, -407, 8130, -2366, -7323, 4870, 5652, -6811, -3310, 7951, 564, -8146, 2257, 7361, -4818, -5684, 6800, 3305, -7958, -514, 8137, -2352, -7308, 4933, 5561, -6906, -3109, 8010, 253, -8101, 2644, 7152, -5212, -5279, 7112, 2712, -8092, 217, 8012, -3128, -6875, 5633, 4817, -7395, -2108, 8167, -895, -7838, 3785, 6438, -6169, -4152, 7709, 1283, -8188, 1771, 7524, -4589, -5804, 6768, 3255, -7996, -238, 8084, -2826, -7013, 5489, 4922, -7366, -2110, 8172, -1022, -7780, 4011, 6234, -6416, -3757, 7868, 707, -8143, 2456, 7185, -5259, -5132, 7265, 2284, -8162, 923, 7797, -3998, -6219, 6456, 3660, -7909, -519, 8114, -2717, -7030, 5526, 4815, -7458, -1820, 8189, -1480, -7592, 4547, 5750, -6879, -2958, 8080, -334, -7944, 3578, 6479, -6234, -3922, 7844, 692, -8130, 2663, 7027, -5573, -4717, 7530, 1583, -8191, 1832, 7423, -4939, -5355, 7184, 2334, -8167, 1107, 7698, -4362, -5853, 6842, 2946, -8095, 499, 7880, -3865, -6228, 6531, 3426, -8003, 15, 7995, -3465, -6499, 6274, 3779, -7914, -342, 8061, -3171, -6679, 6087, 4014, -7847, -572, 8096, -2991, -6779, 5980, 4135, -7811, -676, 8109, -2928, -6807, 5959, 4147, -7812, -653, 8103, -2983, -6764, 6024, 4049, -7851, -504, 8077, -3155, -6647, 6172, 3839, -7920, -228, 8023, -3441, -6448, 6395, 3511, -8010, 175, 7928, -3834, -6156, 6681, 3059, -8101, 703, 7772, -4325, -5756, 7011, 2476, -8171, 1354, 7533, -4897, -5229, 7360, 1754, -8189, 2119, 7183, -5528, -4558, 7694, 893, -8121, 2983, 6693, -6188, -3728, 7975, -106, -7925, 3922, 6031, -6836, -2726, 8154, -1228, -7558, 4900, 5172, -7421, -1552, 8178, -2449, -6979, 5869, 4096, -7883, -217, 7988, -3725, -6149, 6765, 2797, -8152, 1249, 7530, -4997, -5041, 7510, 1288, -8155, 2794, 6752, -6184, -3645, 8016, -395, -7818, 4341, 5621, -7188, -1979, 8190, -2183, -7080, 5787, 4127, -7895, -93, 7941, -3976, -5902, 7005, 2298, -8189, 1921, 7196, -5639, -4280, 7854, 207, -7962, 3929, 5916, -7011, -2261, 8190, -2021, -7132, 5756, 4111, -7916, 49, 7888, -4207, -5669, 7200, 1860, -8185, 2477, 6869, -6127, -3612, 8048, -680, -7686, 4784, 5125, -7529, -1089, 8112, -3271, -6353, 6690, 2745, -8172, 1670, 7267, -5607, -4228, 7900, -66, -7864, 4347, 5492, -7346, -1479, 8153, -2987, -6516, 6562, 2909, -8162, 1585, 7287, -5607, -4189, 7923, -199, -7813, 4533, 5293, -7477, -1131, 8106, -3393, -6211, 6864, 2367, -8191, 2227, 6938, -6129, -3490, 8093, -1076, -7486, 5306, 4482, -7845, -34, 7863, -4435, -5341, 7474, 1078, -8090, 3542, 6062, -7014, -2044, 8184, -2658, -6657, 6487, 2917, -8171, 1798, 7129, -5924, -3699, 8066, -984, -7495, 5341, 4384, -7897, 222, 7765, -4762, -4979, 7677, 476, -7957, 4198, 5486, -7429, -1108, 8081, -3666, -5914, 7164, 1668, -8154, 3171, 6267, -6900, -2160, 8185, -2725, -6558, 6644, 2580, -8190, 2330, 6790, -6411, -2934, 8176, -1994, -6973, 6203, 3221, -8153, 1716, 7111, -6032, -3447, 8126, -1501, -7213, 5898, 3610, -8105, 1346, 7278, -5808, -3716, 8088, -1257, -7315, 5761, 3761, -8083, 1230, 7320, -5761, -3751, 8086, -1269, -7298, 5806, 3681, -8100, 1370, 7243, -5897, -3555, 8121, -1536, -7158, 6029, 3367, -8148, 1762, 7035, -6201, -3119, 8171, -2052, -6872, 6406, 2806, -8189, 2399, 6660, -6641, -2427, 8188, -2804, -6396, 6895, 1978, -8164, 3259) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L21C32_i
    );

    L21C33_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-5500, -7516, 672, 7947, 4422, -5116, -7697, 195, 7822, 4796, -4766, -7833, -218, 7694, 5104, -4457, -7931, -566, 7573, 5353, -4194, -8000, -849, 7465, 5545, -3981, -8047, -1067, 7378, 5686, -3823, -8076, -1220, 7316, 5778, -3720, -8093, -1309, 7281, 5823, -3674, -8099, -1334, 7275, 5823, -3686, -8095, -1295, 7299, 5777, -3756, -8080, -1192, 7351, 5684, -3882, -8053, -1025, 7429, 5543, -4063, -8010, -793, 7530, 5349, -4297, -7946, -496, 7646, 5100, -4580, -7853, -134, 7773, 4790, -4908, -7726, 293, 7900, 4416, -5273, -7553, 784, 8018, 3971, -5667, -7326, 1335, 8115, 3452, -6082, -7034, 1944, 8177, 2855, -6504, -6666, 2603, 8188, 2178, -6918, -6211, 3302, 8131, 1421, -7308, -5659, 4031, 7991, 587, -7654, -5002, 4772, 7748, -318, -7932, -4233, 5506, 7385, -1283, -8120, -3351, 6209, 6887, -2293, -8191, -2358, 6854, 6240, -3325, -8121, -1261, 7409, 5435, -4352, -7883, -76, 7840, 4469, -5340, -7457, 1175, 8112, 3346, -6250, -6823, 2459, 8188, 2079, -7039, -5973, 3738, 8036, 691, -7657, -4904, 4962, 7627, -782, -8057, -3626, 6075, 6942, -2291, -8191, -2166, 7014, 5972, -3778, -8020, -561, 7716, 4726, -5170, -7511, 1129, 8118, 3227, -6389, -6649, 2832, 8162, 1523, -7352, -5439, 4459, 7807, -317, -7977, -3907, 5911, 7028, -2204, -8191, -2108, 7083, 5827, -4028, -7939, -127, 7872, 4237, -5664, -7188, 1924, 8188, 2325, -6984, -5943, 3910, 7962, 198, -7862, -4246, 5679, 7162, -2006, -8191, -2186, 7074, 5797, -4119, -7896, 102, 7948, 3930, -5957, -6947, 2444, 8181, 1681, -7335, -5373, 4635, 7700, -776, -8089, -3271, 6455, 6491, -3222, -8096, -802, 7697, 4619, -5412, -7296, 1807, 8188, 2227, -7093, -5715, 4287, 7816, -460, -8043, -3470, 6350, 6563, -3157, -8099, -775, 7723, 4514, -5542, -7192, 2072, 8190, 1868, -7294, -5369, 4720, 7628, -1074, -8143, -2809, 6805, 6045, -3934, -7913, 185, 8000, 3595, -6305, -6568, 3213, 8078, 579, -7808, -4236, 5827, 6957, -2583, -8161, -1214, 7597, 4738, -5403, -7240, 2057, 8189, 1716, -7400, -5119, 5050, 7433, -1648, -8188, -2091, 7235, 5385, -4787, -7560, 1358, 8175, 2339, -7120, -5551, 4619, 7629, -1193, -8165, -2465, 7062, 5620, -4556, -7651, 1152, 8163, 2469, -7070, -5598, 4596, 7626, -1238, -8171, -2353, 7139, 5480, -4742, -7553, 1446, 8183, 2113, -7267, -5266, 4985, 7422, -1780, -8191, -1749, 7439, 4943, -5320, -7223, 2231, 8175, 1254, -7643, -4505, 5730, 6933, -2796, -8116, -631, 7850, 3934, -6199, -6536, 3460, 7983, -125, -8037, -3223, 6696, 6003, -4208, -7747, 1004, 8161, 2359, -7191, -5316, 5010, 7368, -1997, -8185, -1343, 7638, 4448, -5833, -6814, 3074, 8056, 176, -7987, -3390, 6625, 6046, -4205, -7728, 1119, 8174, 2134, -7327, -5042, 5330, 7149, -2508, -8139, -697, 7865, 3783, -6384, -6281, 3931, 7814, -890, -8161, -2278, 7278, 5093, -5312, -7142, 2562, 8127, 556, -7915, -3584, 6546, 6079, -4233, -7689, 1315, 8187, 1780, -7516, -4614, 5780, 6785, -3236, -7998, 245, 8089, 2768, -7061, -5391, 5062, 7264, -2379, -8143, -620, 7914, 3524, -6625, -5948, 4453, 7570, -1699, -8189, -1271, 7728, 4064, -6263, -6321, 3990, 7752, -1213, -8188, -1711, 7577, 4406, -6014, -6540, 3698, 7846, -932, -8175, -1942, 7494, 4566, -5899, -6626, 3590, 7873, -858, -8172, -1969, 7492, 4550, -5928, -6587, 3669, 7842, -992, -8181, -1793, 7572, 4359, -6098, -6420, 3933, 7743, -1333, -8191, -1409, 7720, 3983, -6396, -6108, 4370, 7554, -1876, -8174, -814, 7906, 3405, -6793, -5625, 4959, 7238, -2610, -8085, -6, 8082, 2609, -7245, -4935, 5663, 6745, -3512, -7865, 1011, 8185, 1579, -7688, -4005, 6427, 6023, -4540, -7444, 2215, 8134, 314, -8038, -2804, 7170, 5016, -5627, -6746, 3558, 7834, -1167, -8191, -1325, 7789, 3683, -6676, -5698, 4961, 7188, -2807, -8029, 410, 8150, 2012, -7555, -4249, 6299, 6105, -4504, -7428, 2328, 8108, 36, -8099, -2388, 7407, 4529, -6101, -6287, 4295, 7517, -2146, -8131, -171, 8082, 2461, -7387, -4547, 6106, 6262, -4351, -7480, 2262, 8110, -9, -8114, -2236, 7496, 4300, -6316, -6032, 4666, 7305, -2678, -8033, 500, 8168, 1702, -7711, -3774, 6699, 5564, -5217, -6952, 3372, 7845, -1301, -8188, -853, 7964, 2936, -7199, -4811, 5949, 6352, -4308, -7464, 2388, 8076, -321, -8159, -1758, 7712, 3712, -6775, -5422, 5410, 6779, -3714, -7707, 1793, 8152, 226, -8098, -2224, 7550, 4076, -6554, -5676, 5171, 6931, -3494, -7777, 1619, 8165, 337, -8086, -2266, 7546, 4055, -6588, -5610, 5268, 6846, -3666, -7703, 1872, 8137, 11, -8136, -1885, 7702, 3648, -6870, -5214, 5685, 6501, -4217, -7452, 2543, 8021, -752, -8190, -1068, 7953, 2824, -7332, -4435, 6360, 5823, -5093, -6930, 3592, 7705, -1935, -8121, 196, 8163, 1539, -7837, -3197, 7163, 4702, -6178, -5994, 4929, 7017, -3477, -7736, 1884, 8122, -224, -8169, -1438, 7877, 3028, -7268, -4489, 6369, 5759, -5224, -6795, 3881, 7559, -2397, -8030, 830, 8190, 757, -8045, -2308, 7601, 3762, -6885, -5072, 5924, 6189, -4760, -7083, 3435, 7723, -2002, -8094, 508, 8187, 991, -8007, -2448, 7563, 3814, -6877, -5049, 5974, 6112, -4890, -6978, 3659, 7620, -2326, -8027, 931, 8187, 480, -8106, -1869, 7786, 3192, -7247, -4416, 6504, 5504, -5587, -6434, 4521, 7178, -3343, -7727, 2082, 8064, -778, -8191, -538, 8104, 1827, -7815, -3063, 7332, 4212, -6676, -5251, 5862, 6154, -4918, -6908, 3864, 7493, -2733, -7906, 1548, 8136, -340, -8187, -867, 8059, 2043, -7763, -3168, 7306, 4216, -6705, -5171, 5971, 6012, -5128, -6730, 4191, 7309, -3185, -7748, 2125, 8036, -1039, -8177, -58, 8168, 1142, -8018, -2198, 7730, 3205, -7315, -4150, 6782, 5015, -6145, -5794, 5415, 6471, -4609, -7044, 3739, 7502, -2824, -7846, 1875, 8071, -911, -8180, -58, 8173, 1014, -8056, -1948, 7831, 2844, -7508, -3695, 7091, 4489, -6592, -5220, 6016, 5878, -5377, -6461, 4681, 6961, -3942, -7379, 3166, 7708, -2366, -7954, 1550, 8111, -729, -8185, -91, 8175, 898, -8088, -1687, 7924, 2449, -7691, -3181, 7390, 3873, -7030, -4524, 6614, 5126, -6151, -5680, 5643, 6180, -5099, -6627, 4523, 7016, -3924, -7350, 3304, 7626, -2672, -7847, 2030, 8010, -1386, -8122, 741, 8180, -105, -8189, -524, 8148, 1138, -8064, -1737, 7935, 2315, -7769, -2873, 7564, 3404, -7328, -3912, 7059, 4390, -6765, -4842, 6444, 5262, -6105, -5654, 5745, 6014, -5372, -6346, 4985, 6645, -4589, -6917, 4184, 7158, -3776, -7372, 3364, 7557, -2952, -7718, 2539, 7851, -2131, -7961, 1726, 8047, -1328, -8113, 935, 8157, -552, -8183, 177, 8190, 187, -8183, -542, 8159, 884, -8124, -1215, 8074, 1533, -8016, -1840, 7946, 2133, -7869, -2414, 7784, 2681, -7694, -2937, 7598, 3179, -7499, -3409, 7396, 3626, -7293, -3831, 7187, 4023, -7082, -4205, 6976, 4374, -6874, -4534, 6771, 4680, -6673, -4818, 6577, 4944, -6485, -5061, 6397, 5167, -6314, -5266, 6235, 5354, -6164, -5435, 6096, 5505, -6036, -5569, 5980, 5622, -5933, -5670, 5891, 5708, -5858, -5741, 5830, 5764, -5811, -5781, 5797, 5789, -5793, -5792, 5793, 5786, -5804, -5774, 5819, 5753, -5844, -5726, 5873, 5690, -5912, -5648, 5956, 5596, -6008, -5538, 6065, 5470, -6129, -5396, 6198, 5311, -6275, -5218, 6354, 5115, -6441, -5004, 6530, 4882, -6625, -4751, 6722, 4608, -6823, -4456, 6925, 4291, -7030, -4116, 7134, 3928, -7240, -3730, 7344, 3518, -7449, -3296, 7548, 3059, -7647, -2811, 7739, 2549, -7828, -2276, 7908, 1987, -7982, -1689, 8046, 1375, -8101, -1051, 8143, 713, -8174, -366, 8188, 6, -8190, 363, 8172, -743, -8138, 1130, 8082, -1527, -8008, 1927, 7908, -2335, -7788, 2745, 7640, -3158, -7469, 3570, 7268, -3982, -7042, 4387, 6784, -4789, -6500, 5180, 6183, -5561, -5838, 5927, 5461, -6278, -5056, 6607, 4619, -6916, -4155, 7197, 3661, -7451, -3142, 7671, 2596, -7858, -2029, 8004, 1439, -8112, -833, 8174, 210, -8191, 422, 8157, -1064, -8073, 1708, 7935, -2352, -7743, 2989, 7494, -3617, -7190, 4226, 6828, -4816, -6411, 5375, 5936, -5903, -5410, 6388, 4830, -6830, -4204, 7217, 3531, -7549, -2819, 7816, 2071, -8016, -1295, 8141, 495, -8191, 318, 8158, -1140, -8043, 1959, 7841, -2769, -7555, 3558, 7180, -4318, -6721, 5035, 6178, -5705, -5558, 6313, 4862, -6852, -4099, 7310, 3275, -7682, -2401, 7956, 1483, -8129, -538, 8190, -427, -8141, 1394, 7973, -2354, -7689, 3287, 7287, -4182, -6772, 5021, 6145, -5791, -5416, 6476, 4592, -7063, -3686, 7538, 2707, -7891, -1675, 8110, 602, -8191, 490, 8124, -1586, -7911, 2660, 7546, -3697, -7037, 4670, 6386, -5564, -5606, 6353, 4705, -7023, -3702, 7554, 2612, -7933, -1460, 8145, 264, -8184, 946, 8043, -2147, -7722, 3307, 7221, -4404, -6551, 5405, 5720, -6288, -4747, 7025, 3649, -7598, -2454, 7984, 1186, -8174, 120, 8153, -1435, -7922, 2720, 7477, -3945, -6830, 5071, 5989, -6067, -4978, 6899, 3817, -7544, -2541, 7975, 1179, -8177, 225, 8137, -1635, -7854, 3003, 7327, -4291, -6572, 5453, 5602, -6452, -4450, 7249, 3144, -7817, -1728, 8130, 242, -8176, 1259, 7942, -2730, -7436, 4115, 6665, -5366, -5656, 6433, 4436, -7277, -3050, 7859, 1540, -8156, 36, 8148, -1621, -7833, 3153, 7212, -4575, -6309, 5825, 5149, -6853, -3778, 7610, 2244, -8065, -611, 8187, -1060, -7972, 2694, 7416, -4226, -6542, 5583, 5377, -6708, -3972, 7541, 2381, -8046, -676, 8188, -1072, -7960, 2779, 7360, -4369, -6415, 5760, 5160, -6888, -3652, 7688, 1958, -8122, -160, 8156, -1658, -7786, 3401, 7021, -4983, -5896, 6318, 4460, -7334, -2786, 7971, 954, -8191, 937, 7973, -2789, -7325, 4497, 6271, -5970, -4867, 7117, 3182, -7872, -1311, 8184, -646, -8030, 2575, 7408, -4365, -6351, 5906, 4912, -7106, -3174, 7883, 1234, -8188, 789, 7991, -2776, -7301, 4598, 6148, -6142, -4604, 7301, 2757, -8001, -725, 8184, -1366, -7835, 3376, 6965, -5173, -5629, 6630, 3906, -7648, -1911, 8146, -226, -8087, 2356, 7464, -4333, -6315, 6012, 4710, -7271, -2764, 8012, 606, -8176, 1603, 7740, -3707, -6732, 5542, 5214, -6973, -3300, 7880, 1123, -8191, 1147, 7871, -3340, -6940, 5280, 5458, -6815, -3540, 7812, 1328, -8190, 997, 7904, -3254, -6974, 5252, 5464, -6826, -3496, 7835, 1224, -8191, 1158, 7852, -3454, -6841, 5461, 5234, -7004, -3166, 7940, 809, -8181, 1627, 7694, -3929, -6517, 5885, 4744, -7317, -2533, 8083, 79, -8108, 2391, 7376, -4649, -5952, 6476, 3957, -7697, -1578, 8185, -963, -7886, 3419, 6817, -5553, -5077, 7146, 2827, -8038, -288, 8128, -2291, -7400, 4647, 5916, -6539, -3822, 7764, 1324, -8191, 1320, 7763, -3836, -6518, 5956, 4576, -7451, -2139, 8150, -539, -7973, 3167, 6926, -5460, -5117, 7158, 2733, -8070, -39, 8081, -2672, -7184, 5088, 5467, -6936, -3121, 7992, 405, -8131, 2365, 7322, -4871, -5653, 6811, 3308, -7952, -564, 8145, -2259, -7362, 4818, 5682, -6802, -3305, 7957, 512, -8138, 2352, 7307, -4935, -5561, 6905, 3107, -8011, -253, 8100, -2646, -7153, 5211, 5277, -7113, -2712, 8092, -218, -8013, 3128, 6873, -5634, -4817, 7395, 2106, -8168, 895, 7837, -3787, -6438, 6168, 4150, -7710, -1283, 8187, -1773, -7525, 4589, 5802, -6770, -3255, 7995, 236, -8085, 2826, 7011, -5491, -4922, 7366, 2108, -8173, 1022, 7779, -4013, -6235, 6416, 3755, -7869, -707, 8142, -2458, -7185, 5259, 5130, -7266, -2284, 8161, -925, -7798, 3998, 6217, -6458, -3660, 7908, 517, -8114, 2717, 7028, -5528, -4815, 7457, 1818, -8190, 1480, 7591, -4549, -5750, 6879, 2956, -8081, 334, 7943, -3580, -6479, 6233, 3920, -7845, -692, 8128, -2665, -7027, 5573, 4715, -7532, -1583, 8190, -1834, -7424, 4939, 5353, -7186, -2334, 8166, -1109, -7699, 4362, 5851, -6843, -2946, 8094, -501, -7881, 3865, 6226, -6533, -3426, 8002, -17, -7995, 3465, 6497, -6276, -3779, 7914, 340, -8062, 3171, 6677, -6089, -4014, 7846, 570, -8097, 2991, 6778, -5982, -4135, 7810, 674, -8110, 2928, 6805, -5961, -4147, 7812, 651, -8104, 2983, 6762, -6026, -4049, 7850, 502, -8078, 3155, 6645, -6174, -3839, 7920, 226, -8024, 3441, 6447, -6397, -3511, 8009, -177, -7928, 3834, 6155, -6683, -3059, 8100, -706, -7773, 4325, 5754, -7013, -2475, 8170, -1357, -7534, 4897, 5227, -7361, -1754, 8188, -2122, -7184, 5528, 4556, -7696, -892, 8119, -2985, -6693, 6188, 3726, -7976, 106, 7923, -3924, -6031, 6835, 2724, -8155, 1228, 7557, -4902, -5172, 7421, 1550, -8178, 2449, 6977, -5871, -4096, 7882, 215, -7989, 3725, 6147, -6766, -2797, 8151, -1251, -7530, 4997, 5039, -7511, -1288, 8153, -2796, -6752, 6184, 3643, -8018, 395, 7816, -4343, -5621, 7187, 1977, -8191, 2184, 7078, -5789, -4127, 7894, 91, -7941, 3976, 5900, -7007, -2298, 8188, -1923, -7196, 5639, 4278, -7855, -207, 7961, -3931, -5916, 7011, 2258, -8191, 2022, 7131, -5758, -4111, 7915, -52, -7889, 4208, 5667, -7202, -1860, 8184, -2479, -6869, 6127, 3609, -8049, 680, 7684, -4787, -5125, 7529, 1087, -8113, 3271, 6351, -6692, -2744, 8171, -1672, -7267, 5607, 4226, -7901, 66, 7863, -4350, -5492, 7346, 1477, -8154, 2987, 6514, -6564, -2908, 8162, -1587, -7287, 5607, 4187, -7924, 199, 7811, -4535, -5293, 7477, 1128, -8106, 3393, 6209, -6866, -2366, 8190, -2229, -6939, 6129, 3488, -8094, 1077, 7484, -5308, -4482, 7845, 32, -7863, 4435, 5338, -7476, -1078, 8089, -3545, -6062, 7014, 2041, -8185, 2658, 6655, -6489, -2917, 8170, -1801, -7129, 5924, 3697, -8068, 984, 7494, -5343, -4384, 7896, -224, -7766, 4763, 4977, -7679, -475, 7956, -4201, -5485, 7429, 1105, -8081, 3666, 5912, -7166, -1667, 8153, -3174, -6267, 6900, 2157, -8186, 2726, 6556, -6646, -2579, 8189, -2333, -6790, 6411, 2932, -8177, 1995, 6971, -6205, -3221, 8152, -1718, -7111, 6032, 3445, -8128, 1501, 7211, -5900, -3610, 8104, -1349, -7278, 5808, 3713, -8089, 1258, 7313, -5763, -3761, 8082, -1233, -7320, 5762, 3749, -8087, 1270, 7296, -5808, -3681, 8100, -1372, -7243, 5897, 3553, -8122, 1536, 7156, -6031, -3367, 8147, -1765, -7035, 6201, 3117, -8172, 2052, 6870, -6408, -2805, 8188, -2401, -6660, 6641, 2425, -8189, 2804, 6394, -6897, -1978, 8163, -3261) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L21C33_i
    );

    L32_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (134, 7798, 4876, -4668, -7873, -381, 7629, 5266, -4259, -7992, -851, 7448, 5606, -3872, -8076, -1275, 7264, 5898, -3513, -8133, -1654, 7083, 6147, -3186, -8167, -1987, 6910, 6357, -2893, -8185, -2275, 6750, 6530, -2636, -8191, -2519, 6607, 6671, -2418, -8190, -2720, 6485, 6782, -2240, -8185, -2878, 6386, 6866, -2102, -8178, -2995, 6312, 6924, -2006, -8172, -3072, 6265, 6959, -1951, -8169, -3108, 6245, 6970, -1938, -8168, -3104, 6254, 6959, -1968, -8171, -3060, 6290, 6924, -2039, -8177, -2976, 6353, 6866, -2151, -8183, -2851, 6442, 6783, -2305, -8189, -2684, 6555, 6672, -2499, -8191, -2475, 6689, 6531, -2732, -8187, -2223, 6843, 6358, -3004, -8172, -1926, 7011, 6149, -3310, -8141, -1585, 7189, 5900, -3651, -8090, -1197, 7373, 5608, -4021, -8012, -764, 7556, 5269, -4417, -7901, -285, 7731, 4879, -4834, -7750, 237, 7890, 4435, -5266, -7551, 802, 8025, 3934, -5705, -7298, 1405, 8125, 3374, -6143, -6984, 2043, 8182, 2753, -6570, -6600, 2709, 8184, 2072, -6975, -6142, 3394, 8119, 1332, -7345, -5604, 4089, 7978, 539, -7667, -4981, 4782, 7748, -304, -7925, -4273, 5459, 7420, -1185, -8103, -3478, 6104, 6984, -2095, -8187, -2600, 6698, 6434, -3018, -8160, -1645, 7221, 5764, -3936, -8007, -622, 7653, 4972, -4830, -7715, 453, 7971, 4062, -5673, -7272, 1563, 8154, 3039, -6441, -6670, 2684, 8181, 1916, -7105, -5907, 3790, 8032, 710, -7636, -4983, 4849, 7692, -555, -8003, -3908, 5826, 7151, -1849, -8180, -2696, 6683, 6402, -3135, -8140, -1371, 7382, 5450, -4373, -7864, 36, 7884, 4304, -5516, -7338, 1484, 8153, 2988, -6516, -6558, 2926, 8159, 1533, -7323, -5530, 4307, 7876, -18, -7888, -4271, 5567, 7293, -1611, -8168, -2814, 6644, 6407, -3182, -8127, -1204, 7477, 5233, -4661, -7742, 498, 8009, 3801, -5971, -7002, 2220, 8190, 2159, -7038, -5918, 3880, 7986, 374, -7788, -4518, 5387, 7378, -1472, -8160, -2853, 6649, 6370, -3282, -8106, -997, 7579, 4991, -4952, -7598, 956, 8100, 3296, -6372, -6637, 2895, 8152, 1368, -7439, -5253, 4698, 7702, -687, -8060, -3507, 6237, 6745, -2738, -8166, -1493, 7393, 5317, -4646, -7717, 663, 8059, 3489, -6264, -6712, 2813, 8157, 1372, -7454, -5192, 4796, 7645, -889, -8100, -3246, 6445, 6529, -3122, -8118, -1005, 7607, 4865, -5141, -7471, 1358, 8158, 2764, -6763, -6178, 3648, 8016, 386, -7822, -4319, 5653, 7155, -2067, -8191, -2034, 7174, 5618, -4370, -7799, 481, 8039, 3519, -6290, -6645, 2991, 8128, 1037, -7616, -4806, 5239, 7394, -1591, -8180, -2441, 6978, 5873, -4092, -7884, 223, 7993, 3692, -6186, -6719, 2903, 8136, 1066, -7617, -4777, 5293, 7349, -1723, -8187, -2248, 7097, 5684, -4349, -7787, 587, 8070, 3303, -6480, -6423, 3391, 8052, 473, -7826, -4225, 5802, 7000, -2457, -8175, -1445, 7486, 5010, -5102, -7438, 1567, 8181, 2313, -7087, -5669, 4404, 7751, -744, -8103, -3077, 6653, 6207, -3735, -7964, -3, 7962, 3733, -6215, -6642, 3110, 8094, 665, -7785, -4291, 5788, 6981, -2546, -8164, -1240, 7589, 4752, -5393, -7245, 2048, 8189, 1725, -7396, -5128, 5039, 7441, -1627, -8188, -2123, 7216, 5421, -4741, -7585, 1283, 8169, 2434, -7064, -5643, 4502, 7684, -1023, -8148, -2662, 6945, 5796, -4332, -7749, 844, 8128, 2807, -6869, -5889, 4230, 7782, -751, -8119, -2874, 6836, 5920, -4202, -7790, 740, 8118, 2860, -6852, -5894, 4245, 7769, -816, -8130, -2768, 6911, 5807, -4361, -7722, 973, 8148, 2593, -7016, -5659, 4545, 7641, -1217, -8171, -2338, 7155, 5443, -4796, -7522, 1540, 8187, 1996, -7327, -5156, 5106, 7352, -1946, -8189, -1569, 7516, 4788, -5469, -7126, 2425, 8160, 1052, -7713, -4334, 5871, 6827, -2976, -8089, -449, 7899, 3785, -6302, -6444, 3587, 7953, -244, -8057, -3137, 6741, 5960, -4249, -7737, 1018, 8161, 2382, -7170, -5365, 4940, 7415, -1867, -8190, -1523, 7559, 4645, -5644, -6972, 2772, 8112, 560, -7883, -3794, 6328, 6384, -3719, -7904, 493, 8105, 2807, -6964, -5638, 4675, 7533, -1624, -8191, -1689, 7509, 4718, -5608, -6978, 2800, 8102, 451, -7923, -3626, 6471, 6212, -3991, -7806, 879, 8155, 2363, -7218, -5229, 5144, 7266, -2270, -8164, -954, 7787, 4021, -6206, -6462, 3667, 7900, -572, -8125, -2607, 7106, 5380, -5010, -7332, 2157, 8170, 1013, -7778, -4027, 6219, 6430, -3737, -7873, 703, 8143, 2427, -7212, -5195, 5221, 7193, -2471, -8138, -634, 7896, 3640, -6512, -6115, 4191, 7703, -1275, -8187, -1819, 7500, 4646, -5751, -6810, 3192, 8008, -190, -8080, -2833, 7021, 5454, -4988, -7312, 2267, 8155, 759, -7874, -3676, 6514, 6083, -4269, -7658, 1448, 8190, 1560, -7619, -4355, 6023, 6557, -3628, -7883, 754, 8157, 2212, -7354, -4882, 5584, 6903, -3088, -8020, 194, 8089, 2718, -7113, -5273, 5221, 7144, -2665, -8097, -227, 8016, 3082, -6920, -5543, 4952, 7298, -2368, -8137, -508, 7957, 3312, -6792, -5702, 4788, 7381, -2202, -8154, -649, 7926, 3413, -6739, -5758, 4737, 7402, -2171, -8155, -650, 7930, 3385, -6764, -5715, 4799, 7362, -2275, -8143, -511, 7967, 3230, -6867, -5569, 4973, 7257, -2512, -8110, -233, 8030, 2943, -7039, -5314, 5252, 7077, -2879, -8043, 186, 8105, 2518, -7266, -4939, 5623, 6806, -3367, -7922, 744, 8168, 1950, -7526, -4429, 6069, 6421, -3964, -7721, 1437, 8190, 1234, -7789, -3770, 6562, 5900, -4650, -7407, 2254, 8135, 369, -8017, -2949, 7069, 5217, -5398, -6945, 3177, 7959, -641, -8164, -1956, 7543, 4348, -6167, -6299, 4176, 7616, -1778, -8176, -793, 7927, 3276, -6903, -5435, 5206, 7057, -3010, -7994, 527, 8157, 1997, -7540, -4327, 6205, 6237, -4288, -7555, 1970, 8158, 525, -7999, -2966, 7095, 5123, -5539, -6805, 3477, 7856, -1104, -8190, -1364, 7779, 3701, -6670, -5701, 4964, 7183, -2821, -8025, 433, 8153, 1985, -7566, -4225, 6317, 6088, -4524, -7420, 2344, 8107, 30, -8099, -2397, 7399, 4552, -6076, -6317, 4243, 7546, -2062, -8142, -287, 8059, 2603, -7313, -4700, 5967, 6405, -4140, -7586, 1980, 8148, 331, -8055, -2611, 7317, 4675, -6001, -6364, 4213, 7544, -2102, -8133, -169, 8085, 2419, -7414, -4477, 6173, 6184, -4466, -7417, 2422, 8083, -204, -8140, -2025, 7586, 4094, -6471, -5856, 4880, 7179, -2937, -7974, 783, 8184, 1418, -7804, -3513, 6862, 5348, -5435, -6798, 3625, 7761, -1567, -8177, -597, 8019, 2711, -7306, -4632, 6090, 6227, -4462, -7393, 2533, 8052, -441, -8168, -1676, 7734, 3672, -6788, -5421, 5394, 6804, -3652, -7739, 1675, 8165, 402, -8064, -2448, 7444, 4329, -6352, -5931, 4860, 7150, -3068, -7919, 1088, 8190, 950, -7955, -2926, 7229, 4713, -6067, -6210, 4538, 7324, -2742, -7996, 787, 8188, 1207, -7895, -3124, 7138, 4850, -5967, -6290, 4453, 7359, -2689, -8004, 775, 8188, 1174, -7910, -3052, 7187, 4750, -6066, -6181, 4612, 7263, -2911, -7945, 1054, 8190, 850, -7993, -2705, 7367, 4406, -6352, -5869, 5003, 7015, -3398, -7793, 1620, 8161, 234, -8109, -2071, 7640, 3793, -6787, -5320, 5593, 6571, -4126, -7492, 2457, 8038, -675, -8188, -1135, 7937, 2881, -7305, -4484, 6323, 5864, -5046, -6963, 3533, 7728, -1862, -8131, 109, 8154, 1641, -7804, -3310, 7097, 4821, -6073, -6110, 4778, 7119, -3278, -7810, 1637, 8153, 68, -8139, -1765, 7772, 3377, -7074, -4840, 6075, 6089, -4825, -7079, 3376, 7768, -1794, -8134, 143, 8162, 1505, -7859, -3088, 7238, 4537, -6332, -5802, 5176, 6830, -3823, -7587, 2324, 8044, -743, -8191, -861, 8022, 2424, -7552, -3891, 6798, 5203, -5795, -6319, 4581, 7196, -3207, -7809, 1720, 8135, -180, -8170, -1362, 7913, 2847, -7380, -4228, 6591, 5454, -5580, -6488, 4379, 7295, -3038, -7854, 1599, 8145, -115, -8167, -1368, 7919, 2798, -7416, -4132, 6674, 5325, -5724, -6346, 4596, 7160, -3330, -7748, 1966, 8093, -549, -8190, -880, 8036, 2273, -7644, -3593, 7024, 4799, -6203, -5861, 5202, 6745, -4059, -7433, 2803, 7904, -1476, -8153, 112, 8171, 1246, -7965, -2565, 7541, 3806, -6917, -4940, 6109, 5935, -5145, -6770, 4049, 7422, -2856, -7882, 1594, 8135, -300, -8184, -997, 8026, 2260, -7672, -3463, 7130, 4573, -6421, -5569, 5559, 6425, -4572, -7127, 3482, 7657, -2319, -8009, 1107, 8176, 121, -8159, -1342, 7958, 2524, -7585, -3646, 7046, 4681, -6361, -5611, 5543, 6416, -4615, -7083, 3593, 7599, -2506, -7958, 1373, 8152, -220, -8184, -932, 8052, 2057, -7767, -3137, 7331, 4149, -6761, -5078, 6065, 5905, -5263, -6619, 4367, 7207, -3400, -7663, 2376, 7979, -1318, -8154, 242, 8185, 829, -8078, -1881, 7833, 2893, -7462, -3852, 6967, 4740, -6366, -5548, 5664, 6261, -4879, -6872, 4022, 7371, -3110, -7755, 2155, 8019, -1177, -8163, 186, 8185, 799, -8090, -1767, 7878, 2702, -7560, -3594, 7137, 4429, -6621, -5200, 6018, 5893, -5341, -6506, 4598, 7028, -3803, -7458, 2964, 7789, -2095, -8023, 1206, 8155, -310, -8190, -584, 8126, 1462, -7969, -2319, 7721, 3141, -7388, -3922, 6975, 4653, -6490, -5329, 5937, 5940, -5328, -6486, 4666, 6959, -3963, -7359, 3225, 7680, -2463, -7925, 1681, 8089, -892, -8177, 99, 8185, 686, -8121, -1459, 7982, 2211, -7775, -2939, 7501, 3632, -7167, -4291, 6774, 4906, -6331, -5478, 5839, 5998, -5307, -6468, 4737, 6882, -4138, -7242, 3512, 7543, -2869, -7788, 2209, 7973, -1542, -8102, 869, 8173, -200, -8190, -467, 8152, 1121, -8063, -1764, 7923, 2386, -7737, -2990, 7505, 3567, -7232, -4119, 6919, 4639, -6573, -5129, 6192, 5585, -5784, -6007, 5349, 6391, -4892, -6740, 4415, 7049, -3924, -7322, 3418, 7556, -2904, -7753, 2381, 7912, -1856, -8035, 1327, 8121, -802, -8174, 279, 8190, 237, -8177, -747, 8130, 1245, -8055, -1734, 7949, 2208, -7819, -2669, 7663, 3113, -7484, -3542, 7282, 3951, -7062, -4344, 6822, 4716, -6567, -5071, 6296, 5403, -6013, -5718, 5716, 6010, -5411, -6284, 5096, 6536, -4776, -6769, 4448, 6982, -4117, -7176, 3781, 7350, -3446, -7508, 3107, 7645, -2771, -7767, 2434, 7870, -2101, -7960, 1769, 8032, -1443, -8091, 1120, 8134, -803, -8166, 490, 8184, -185, -8191, -115, 8186, 406, -8173, -691, 8148, 967, -8117, -1237, 8075, 1497, -8029, -1750, 7973, 1993, -7914, -2230, 7848, 2456, -7779, -2675, 7704, 2884, -7628, -3086, 7547, 3278, -7465, -3463, 7380, 3638, -7296, -3807, 7209, 3966, -7124, -4119, 7037, 4262, -6952, -4399, 6867, 4527, -6785, -4650, 6702, 4764, -6624, -4872, 6546, 4972, -6472, -5067, 6400, 5154, -6332, -5237, 6266, 5311, -6205, -5382, 6146, 5444, -6093, -5503, 6042, 5554, -5998, -5602, 5955, 5643, -5919, -5680, 5886, 5710, -5859, -5737, 5835, 5757, -5818, -5774, 5804, 5784, -5796, -5791, 5792, 5791, -5794, -5789, 5799, 5779, -5811, -5767, 5826, 5747, -5847, -5725, 5872, 5695, -5903, -5662, 5936, 5623, -5977, -5579, 6019, 5529, -6068, -5475, 6119, 5413, -6176, -5348, 6235, 5274, -6299, -5197, 6365, 5111, -6436, -5021, 6508, 4923, -6585, -4819, 6662, 4707, -6744, -4590, 6825, 4464, -6910, -4332, 6994, 4191, -7081, -4044, 7166, 3887, -7253, -3724, 7338, 3551, -7424, -3372, 7506, 3183, -7588, -2987, 7666, 2780, -7742, -2567, 7814, 2343, -7882, -2113, 7944, 1872, -8002, -1625, 8052, 1368, -8098, -1104, 8133, 830, -8162, -550, 8180, 261, -8191, 34, 8188, -337, -8177, 645, 8151, -961, -8115, 1280, 8062, -1606, -7998, 1934, 7917, -2268, -7821, 2602, 7708, -2940, -7579, 3276, 7431, -3614, -7266, 3949, 7081, -4283, -6878, 4612, 6655, -4937, -6413, 5254, 6149, -5565, -5867, 5865, 5563, -6156, -5240, 6433, 4896, -6697, -4533, 6944, 4150, -7175, -3750, 7385, 3329, -7577, -2894, 7744, 2440, -7888, -1973, 8005, 1491, -8096, -998, 8156, 493, -8188, 19, 8186, -540, -8152, 1064, 8082, -1592, -7979, 2118, 7837, -2643, -7660, 3161, 7443, -3673, -7191, 4171, 6898, -4656, -6570, 5123, 6203, -5570, -5801, 5991, 5361, -6387, -4889, 6750, 4382, -7081, -3847, 7373, 3281, -7627, -2691, 7835, 2077, -8000, -1445, 8113, 795, -8178, -135, 8188, -535, -8145, 1205, 8044, -1877, -7888, 2540, 7672, -3193, -7400, 3828, 7069, -4442, -6682, 5026, 6239, -5578, -5745, 6090, 5197, -6559, -4605, 6977, 3966, -7342, -3290, 7645, 2578, -7887, -1838, 8060, 1074, -8163, -295, 8190, -496, -8143, 1287, 8016, -2074, -7813, 2846, 7529, -3598, -7169, 4319, 6731, -5003, -6223, 5639, 5642, -6222, -4999, 6740, 4294, -7192, -3538, 7564, 2734, -7857, -1895, 8059, 1025, -8171, -138, 8185, -759, -8102, 1652, 7918, -2533, -7636, 3387, 7254, -4207, -6779, 4977, 6210, -5689, -5557, 6329, 4823, -6891, -4020, 7360, 3154, -7733, -2240, 7998, 1286, -8152, -308, 8188, -682, -8107, 1668, 7902, -2637, -7578, 3571, 7135, -4459, -6580, 5281, 5916, -6027, -5156, 6679, 4305, -7229, -3381, 7663, 2392, -7973, -1359, 8148, 294, -8188, 781, 8084, -1851, -7839, 2893, 7452, -3892, -6930, 4825, 6277, -5677, -5505, 6427, 4625, -7063, -3653, 7566, 2604, -7929, -1499, 8137, 357, -8189, 797, 8075, -1944, -7799, 3056, 7360, -4114, -6768, 5091, 6030, -5968, -5161, 6721, 4175, -7336, -3095, 7792, 1938, -8081, -735, 8190, -494, -8116, 1717, 7856, -2909, -7414, 4038, 6796, -5081, -6016, 6007, 5086, -6796, -4031, 7423, 2870, -7873, -1635, 8130, 350, -8186, 949, 8034, -2232, -7678, 3463, 7119, -4612, -6374, 5644, 5456, -6534, -4389, 7252, 3197, -7780, -1914, 8095, 570, -8191, 795, 8057, -2146, -7697, 3442, 7115, -4647, -6327, 5722, 5350, -6638, -4213, 7360, 2944, -7870, -1584, 8143, 166, -8173, 1261, 7951, -2658, -7484, 3977, 6780, -5180, -5860, 6223, 4748, -7073, -3480, 7698, 2092, -8076, -631, 8190, -860, -8034, 2327, 7606, -3724, -6922, 5000, 5997, -6112, -4863, 7015, 3553, -7681, -2115, 8077, 594, -8190, 953, 8008, -2474, -7538, 3911, 6789, -5212, -5789, 6325, 4569, -7209, -3173, 7823, 1651, -8146, -60, 8157, -1541, -7855, 3087, 7244, -4522, -6348, 5782, 5196, -6820, -3833, 7586, 2309, -8052, -686, 8189, -973, -7993, 2597, 7462, -4122, -6620, 5478, 5494, -6609, -4131, 7462, 2585, -7999, -923, 8190, -789, -8026, 2470, 7506, -4051, -6653, 5455, 5497, -6622, -4090, 7492, 2490, -8025, -772, 8190, -991, -7977, 2712, 7389, -4315, -6453, 5718, 5205, -6856, -3706, 7667, 2021, -8113, -233, 8163, -1575, -7814, 3311, 7076, -4890, -5984, 6228, 4586, -7260, -2952, 7925, 1160, -8188, 696, 8029, -2525, -7454, 4227, 6485, -5715, -5173, 6904, 3579, -7732, -1791, 8146, -102, -8123, 1995, 7656, -3787, -6769, 5375, 5504, -6673, -3930, 7601, 2128, -8107, -202, 8154, -1744, -7738, 3596, 6874, -5248, -5612, 6600, 4017, -7572, -2183, 8101, 212, -8154, 1777, 7718, -3667, -6819, 5342, 5504, -6699, -3850, 7650, 1954, -8136, 68, 8118, -2094, -7595, 3994, 6593, -5651, -5172, 6953, 3416, -7817, -1438, 8181, -642, -8018, 2684, 7331, -4560, -6164, 6141, 4585, -7322, -2698, 8017, 623, -8180, 1498, 7789, -3527, -6870, 5320, 5477, -6756, -3705, 7729, 1669, -8170, 488, 8039, -2619, -7345, 4570, 6128, -6204, -4472, 7399, 2489, -8068, -322, 8153, -1877, -7647, 3943, 6578, -5728, -5023, 7094, 3089, -7937, -920, 8188, -1325, -7825, 3476, 6866, -5371, -5384, 6859, 3482, -7826, -1308, 8189, -976, -7917, 3188, 7023, -5158, -5576, 6725, 3680, -7764, -1488, 8184, -832, -7949, 3090, 7068, -5105, -5612, 6708, 3690, -7767, -1461, 8186, -897, -7928, 3185, 7005, -5215, -5494, 6809, 3512, -7833, -1228, 8190, -1169, -7849, 3470, 6828, -5480, -5214, 7017, 3140, -7947, -786, 8179, -1645, -7690, 3935, 6515, -5883, -4756, 7306, 2562, -8077, -133, 8116, -2317, -7417, 4559, 6034, -6391, -4093, 7635, 1766, -8175, 730, 7950, -3166, -6980, 5308, 5346, -6956, -3202, 7943, 744, -8174, 1789, 7618, -4158, -6324, 6128, 4410, -7508, -2061, 8152, -498, -7996, 3013, 7046, -5237, -5392, 6941, 3193, -7955, -668, 8165, -1933, -7550, 4342, 6161, -6315, -4138, 7641, 1681, -8183, 954, 7874, -3498, -6744, 5681, 4901, -7272, -2538, 8097, -102, -8064, 2736, 7168, -5085, -5501, 6890, 3234, -7956, -613, 8157, -2084, -7468, 4557, 5955, -6536, -3782, 7794, 1183, -8189, 1553, 7668, -4123, -6286, 6233, 4188, -7645, -1612, 8187, -1156, -7797, 3796, 6508, -6008, -4466, 7527, 1899, -8176, 894, 7868, -3590, -6638, 5868, 4619, -7459, -2050, 8165, -772, -7899, 3506, 6682, -5826, -4658, 7445, 2063, -8166, 788, 7889, -3550, -6646, 5880, 4579, -7492, -1942, 8175, -944, -7842, 3717, 6524, -6032, -4384, 7588, 1682, -8188, 1237, 7745, -4007, -6312, 6268, 4062, -7727, -1284, 8188, -1668, -7587, 4408, 5992, -6578, -3608, 7886, 742, -8157, 2227, 7343, -4908, -5551, 6937, 3009, -8041, -58, 8061, -2908, -6991, 5485, 4965, -7320, -2258, 8155, -767, -7871, 3691, 6497, -6112, -4219, 7685, 1346, -8189, 1720, 7543, -4552, -5833, 6745, 3292, -7987, -278, 8091, -2783, -7038, 5450, 4968, -7338, -2178, 8166, -935, -7810, 3917, 6310, -6334, -3884, 7823, 879, -8161, 2261, 7288, -5074, -5330, 7132, 2569, -8129, 582, 7901, -3653, -6481, 6176, 4072, -7766, -1039, 8171, -2161, -7324, 5033, 5346, -7136, -2539, 8135, -671, -7871, 3781, 6373, -6306, -3874, 7842, 757, -8144, 2484, 7153, -5338, -5022, 7344, 2081, -8179, 1198, 7697, -4292, -5971, 6695, 3271, -8016, -35, 8028, -3216, -6726, 5942, 4312, -7696, -1183, 8176, -2151, -7299, 5131, 5199, -7260, -2226, 8171, -1130, -7708, 4299, 5936, -6747, -3153, 8048, -175, -7976, 3478, 6533, -6190, -3962, 7836, 698, -8128, 2691, 7003, -5619, -4653, 7566, 1480, -8188, 1958, 7363, -5058, -5233, 7263, 2166, -8179, 1292, 7631, -4526, -5712, 6950, 2757, -8124, 701, 7823, -4040, -6099, 6645, 3254, -8040, 191, 7956, -3610, -6405, 6365, 3662, -7945, -235, 8044, -3245, -6641, 6120, 3985, -7851, -575, 8100, -2951, -6815, 5922, 4228, -7770, -831, 8132, -2733, -6934, 5776, 4395, -7710, -1002, 8150, -2594, -7006, 5688, 4488, -7676, -1088, 8157, -2534, -7032, 5660, 4511, -7671, -1091, 8156, -2555, -7014, 5693, 4462, -7695, -1009, 8147, -2656, -6952, 5786, 4342, -7747, -843, 8126, -2836, -6843, 5937, 4147, -7821, -592, 8089, -3093, -6680, 6140, 3875, -7912, -256, 8027, -3424, -6458, 6387, 3521, -8008, 165, 7930, -3823, -6166, 6671, 3080, -8097, 670, 7785, -4284, -5796, 6977, 2548, -8164, 1256, 7577, -4795, -5337, 7290, 1922, -8191, 1918, 7289, -5344, -4777, 7591, 1200, -8158, 2648, 6905, -5913, -4109, 7857, 384, -8040, 3432, 6408, -6480, -3325, 8062, -521, -7814, 4252, 5780, -7018, -2421, 8177, -1502, -7456, 5084, 5010, -7496, -1400, 8169, -2543, -6942, 5897, 4088, -7877, -272, 8007, -3616, -6252, 6654, 3012, -8122, 946, 7659, -4686, -5370, 7311, 1790, -8188, 2224, 7095, -5710, -4290, 7819, 439, -8036, 3523, 6295, -6634, -3017, 8125, -1008, -7626, 4789, 5246, -7397, -1569, 8176, -2504, -6929, 5960, 3951, -7935, 16, 7925, -3987, -5927, 6960, 2431, -8182, 1684, 7333, -5379, -4622, 7710, 727, -8078, 3358, 6376, -6590, -3036, 8129, -1094, -7573, 4945, 5054, -7521, -1220, 8142, -2940, -6640, 6335, 3395, -8076, 744, 7692, -4696, -5279, 7410, 1463, -8165, 2746, 6746, -6231, -3526, 8053, -644, -7720, 4646, 5308, -7403, -1462, 8162, -2788, -6710, 6285, 3429, -8076, 790, 7662, -4801, -5148, 7498, 1213, -8135, 3060, 6525, -6495, -3105, 8130, -1184, -7505, 5148, 4782, -7679, -718, 8057, -3557, -6171, 6832, 2538, -8183, 1817, 7213, -5664, -4192, 7901, -31, -7885, 4250, 5607, -7256, -1716, 8175, -2678, -6737, 6301, 3343, -8103, 1026, 7547, -5103, -4790, 7692, 625, -8032, 3727, 6008, -6990, -2211, 8190, -2247, -6968, 6042, 3671, -8047, 723, 7650, -4908, -4964, 7626, 782, -8056, 3639, 6055, -6969, -2221, 8190, -2293, -6927, 6114, 3549, -8076, 917, 7567, -5109, -4736, 7734, 441, -7980, 3994, 5757, -7199, -1747, 8172, -2813, -6602, 6501, 2965, -8161, 1603, 7261, -5676, -4077, 7963, -400, -7739, 4754, 5060, -7607, -771, 8040, -3771, -5909, 7112, 1882, -8179, 2753, 6616, -6509, -2919, 8167, -1728, -7184, 5819, 3865, -8025, 715, 7614, -5069, -4715, 7767, 264, -7919, 4278, 5461, -7417, -1198, 8104, -3469, -6107, 6988, 2073, -8186, 2655, 6649, -6503, -2885, 8173, -1855, -7097, 5974, 3625, -8082, 1076, 7454, -5420, -4295, 7924, -333, -7731, 4851, 4891, -7715, -373, 7931, -4282, -5419, 7463, 1030, -8070, 3719, 5877, -7185, -1640, 8151, -3175, -6275, 6885, 2198, -8188, 2654, 6612, -6579, -2706, 8186, -2163, -6899, 6270, 3161, -8156, 1705, 7136, -5970, -3567, 8103, -1285, -7333, 5681, 3924, -8037, 903, 7492, -5411, -4235, 7961, -565, -7621, 5163, 4501, -7884, 266, 7721, -4943, -4727, 7808, -12, -7801, 4751, 4911, -7739, -200, 7860, -4592, -5059, 7679, 368, -7904, 4465, 5170, -7632, -494, 7933, -4375, -5247, 7598, 574, -7952, 4319, 5289, -7581, -614, 7958, -4302, -5300, 7578, 609, -7956, 4320, 5276, -7594, -562, 7941, -4376, -5220, 7623, 470, -7917, 4466, 5128, -7669, -337, 7878, -4593, -5004, 7726, 159, -7827, 4752, 4840, -7795, 61, 7755, -4945, -4640, 7868, -325, -7664, 5165, 4398, -7947, 631, 7546, -5413, -4114, 8022, -980, -7400, 5683, 3784, -8092, 1369, 7218, -5972, -3408, 8146, -1798, -6998, 6273, 2981, -8183, 2262, 6730, -6582, -2505) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L32_i
    );

    L32C31_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-132, -7798, -4879, 4665, 7873, 382, -7629, -5269, 4256, 7991, 852, -7448, -5609, 3869, 8076, 1277, -7264, -5901, 3510, 8132, 1655, -7082, -6150, 3183, 8166, 1988, -6909, -6359, 2889, 8184, 2276, -6749, -6533, 2633, 8190, 2520, -6607, -6673, 2415, 8189, 2721, -6484, -6784, 2237, 8183, 2880, -6385, -6868, 2099, 8177, 2997, -6311, -6926, 2002, 8171, 3073, -6264, -6961, 1948, 8168, 3109, -6245, -6972, 1935, 8167, 3105, -6253, -6961, 1964, 8170, 3062, -6289, -6927, 2035, 8175, 2977, -6352, -6869, 2148, 8182, 2852, -6441, -6785, 2302, 8188, 2686, -6554, -6674, 2496, 8190, 2477, -6689, -6534, 2729, 8186, 2224, -6842, -6361, 3000, 8171, 1928, -7010, -6152, 3307, 8141, 1586, -7189, -5903, 3647, 8089, 1199, -7373, -5611, 4018, 8012, 765, -7556, -5272, 4414, 7900, 287, -7731, -4882, 4831, 7749, -236, -7890, -4438, 5263, 7551, -801, -8025, -3937, 5702, 7298, -1404, -8126, -3377, 6141, 6984, -2042, -8183, -2756, 6568, 6601, -2707, -8185, -2075, 6973, 6143, -3393, -8121, -1336, 7343, 5605, -4088, -7979, -542, 7665, 4982, -4781, -7750, 300, 7923, 4274, -5459, -7422, 1182, 8102, 3479, -6103, -6986, 2092, 8186, 2601, -6697, -6436, 3015, 8159, 1646, -7221, -5766, 3933, 8007, 624, -7653, -4975, 4827, 7715, -451, -7972, -4065, 5671, 7272, -1561, -8155, -3042, 6439, 6671, -2683, -8182, -1919, 7103, 5908, -3789, -8033, -713, 7634, 4984, -4848, -7694, 552, 8002, 3909, -5825, -7153, 1845, 8178, 2697, -6683, -6405, 3132, 8139, 1372, -7382, -5452, 4370, 7864, -35, -7884, -4307, 5514, 7338, -1483, -8154, -2991, 6514, 6559, -2925, -8160, -1536, 7321, 5531, -4306, -7878, 15, 7886, 4272, -5566, -7295, 1608, 8166, 2815, -6644, -6410, 3179, 8126, 1205, -7477, -5236, 4658, 7741, -497, -8009, -3804, 5969, 7003, -2219, -8191, -2162, 7036, 5918, -3879, -7988, -377, 7787, 4519, -5386, -7380, 1469, 8159, 2854, -6649, -6373, 3279, 8105, 998, -7580, -4994, 4949, 7598, -955, -8101, -3299, 6370, 6638, -2894, -8153, -1371, 7437, 5253, -4697, -7703, 683, 8059, 3507, -6237, -6747, 2735, 8165, 1494, -7393, -5319, 4643, 7717, -662, -8059, -3492, 6262, 6712, -2812, -8158, -1375, 7453, 5193, -4795, -7647, 886, 8099, 3247, -6445, -6531, 3119, 8117, 1006, -7608, -4868, 5139, 7471, -1357, -8159, -2767, 6761, 6178, -3647, -8017, -389, 7821, 4319, -5653, -7157, 2064, 8190, 2035, -7174, -5621, 4367, 7799, -480, -8039, -3521, 6288, 6645, -2990, -8130, -1040, 7614, 4807, -5239, -7396, 1588, 8179, 2442, -6978, -5875, 4089, 7883, -222, -7993, -3695, 6184, 6719, -2902, -8137, -1069, 7616, 4777, -5292, -7351, 1720, 8186, 2249, -7097, -5686, 4346, 7787, -586, -8071, -3305, 6478, 6423, -3390, -8053, -476, 7824, 4225, -5802, -7002, 2454, 8174, 1446, -7486, -5013, 5099, 7438, -1566, -8182, -2315, 7085, 5670, -4403, -7752, 742, 8102, 3077, -6653, -6210, 3733, 7963, 4, -7962, -3736, 6213, 6642, -3110, -8095, -668, 7783, 4292, -5787, -6983, 2543, 8163, 1241, -7589, -4755, 5390, 7245, -2047, -8190, -1728, 7394, 5128, -5039, -7443, 1624, 8186, 2124, -7216, -5423, 4739, 7585, -1282, -8170, -2437, 7062, 5644, -4502, -7686, 1020, 8147, 2663, -6945, -5799, 4330, 7749, -843, -8129, -2810, 6867, 5889, -4230, -7784, 748, 8117, 2875, -6836, -5922, 4199, 7789, -739, -8119, -2862, 6850, 5894, -4244, -7771, 813, 8129, 2768, -6911, -5809, 4358, 7722, -973, -8149, -2595, 7014, 5659, -4544, -7642, 1214, 8170, 2338, -7155, -5445, 4794, 7521, -1539, -8188, -1998, 7325, 5156, -5105, -7354, 1943, 8188, 1570, -7516, -4790, 5466, 7126, -2424, -8162, -1055, 7712, 4335, -5871, -6828, 2974, 8088, 449, -7899, -3788, 6300, 6444, -3587, -7954, 242, 8055, 3138, -6741, -5962, 4246, 7736, -1017, -8162, -2385, 7168, 5365, -4940, -7417, 1864, 8189, 1524, -7560, -4647, 5642, 6972, -2772, -8114, -563, 7882, 3795, -6328, -6386, 3717, 7904, -493, -8105, -2809, 6962, 5638, -4674, -7535, 1621, 8190, 1690, -7509, -4721, 5606, 6977, -2800, -8104, -454, 7921, 3626, -6471, -6214, 3989, 7805, -879, -8156, -2366, 7216, 5229, -5144, -7267, 2268, 8163, 954, -7788, -4024, 6204, 6462, -3667, -7902, 569, 8124, 2607, -7107, -5382, 5008, 7332, -2157, -8171, -1016, 7777, 4027, -6219, -6432, 3735, 7872, -703, -8144, -2429, 7211, 5195, -5221, -7195, 2469, 8137, 635, -7896, -3642, 6511, 6115, -4191, -7705, 1273, 8186, 1819, -7500, -4648, 5749, 6810, -3191, -8009, 188, 8079, 2834, -7021, -5456, 4986, 7312, -2267, -8156, -761, 7873, 3677, -6514, -6085, 4267, 7657, -1448, -8191, -1563, 7617, 4355, -6023, -6559, 3626, 7882, -753, -8158, -2215, 7352, 4882, -5584, -6905, 3086, 8019, -193, -8090, -2720, 7111, 5274, -5221, -7145, 2663, 8097, 228, -8017, -3085, 6918, 5543, -4952, -7300, 2365, 8136, 509, -7958, -3315, 6790, 5702, -4788, -7383, 2200, 8153, 649, -7927, -3415, 6737, 5758, -4737, -7404, 2169, 8154, 650, -7931, -3388, 6763, 5715, -4799, -7364, 2273, 8142, 512, -7968, -3232, 6866, 5569, -4973, -7259, 2510, 8109, 233, -8031, -2945, 7038, 5314, -5252, -7079, 2876, 8042, -186, -8105, -2520, 7265, 4939, -5623, -6807, 3364, 7921, -744, -8168, -1953, 7524, 4429, -6069, -6423, 3962, 7720, -1437, -8191, -1237, 7787, 3771, -6563, -5902, 4648, 7407, -2254, -8136, -371, 8016, 2949, -7069, -5219, 5396, 6945, -3177, -7960, 638, 8163, 1956, -7543, -4350, 6165, 6299, -4176, -7617, 1775, 8175, 793, -7928, -3278, 6901, 5435, -5206, -7058, 3008, 7993, -527, -8157, -2000, 7539, 4327, -6205, -6239, 4286, 7555, -1970, -8159, -527, 7997, 2966, -7095, -5125, 5537, 6805, -3477, -7858, 1102, 8189, 1365, -7780, -3703, 6668, 5700, -4964, -7185, 2819, 8024, -433, -8154, -1988, 7564, 4225, -6317, -6090, 4522, 7419, -2343, -8108, -33, 8098, 2397, -7400, -4554, 6075, 6317, -4243, -7547, 2060, 8141, 287, -8060, -2605, 7311, 4700, -5967, -6407, 4138, 7586, -1980, -8149, -334, 8054, 2611, -7317, -4677, 6000, 6363, -4214, -7546, 2100, 8132, 169, -8086, -2421, 7413, 4477, -6173, -6186, 4464, 7417, -2422, -8084, 202, 8139, 2025, -7586, -4096, 6469, 5855, -4880, -7180, 2935, 7973, -783, -8185, -1420, 7803, 3513, -6863, -5350, 5434, 6798, -3625, -7762, 1565, 8176, 597, -8019, -2713, 7305, 4632, -6090, -6229, 4460, 7393, -2533, -8053, 439, 8167, 1676, -7734, -3674, 6786, 5420, -5394, -6805, 3650, 7738, -1675, -8166, -404, 8063, 2448, -7444, -4331, 6351, 5930, -4860, -7152, 3066, 7919, -1088, -8191, -952, 7954, 2926, -7230, -4715, 6065, 6209, -4538, -7325, 2740, 7996, -787, -8189, -1209, 7894, 3124, -7138, -4852, 5966, 6289, -4453, -7360, 2687, 8003, -776, -8189, -1176, 7909, 3051, -7187, -4752, 6065, 6180, -4612, -7264, 2909, 7944, -1055, -8191, -852, 7992, 2705, -7367, -4407, 6350, 5868, -5003, -7017, 3396, 7792, -1620, -8162, -236, 8108, 2071, -7641, -3795, 6786, 5319, -5594, -6573, 4124, 7492, -2457, -8039, 673, 8187, 1135, -7938, -2883, 7304, 4484, -6324, -5866, 5044, 6963, -3533, -7730, 1860, 8131, -109, -8155, -1643, 7802, 3310, -7097, -4823, 6071, 6110, -4779, -7121, 3276, 7809, -1637, -8154, -70, 8138, 1764, -7773, -3378, 7072, 4839, -6075, -6091, 4823, 7079, -3376, -7769, 1792, 8133, -143, -8163, -1507, 7858, 3088, -7239, -4539, 6331, 5802, -5176, -6831, 3821, 7587, -2324, -8046, 742, 8190, 861, -8023, -2426, 7551, 3890, -6798, -5205, 5794, 6319, -4582, -7198, 3205, 7808, -1720, -8136, 178, 8169, 1362, -7914, -2849, 7379, 4227, -6592, -5455, 5578, 6488, -4380, -7296, 3037, 7853, -1599, -8146, 113, 8166, 1368, -7920, -2799, 7414, 4132, -6674, -5327, 5722, 6345, -4596, -7161, 3329, 7748, -1966, -8094, 547, 8189, 879, -8037, -2274, 7643, 3593, -7025, -4801, 6201, 5860, -5203, -6746, 4057, 7432, -2803, -7906, 1474, 8152, -112, -8172, -1248, 7964, 2565, -7541, -3808, 6915, 4940, -6109, -5936, 5143, 6769, -4050, -7424, 2855, 7881, -1595, -8136, 298, 8183, 996, -8027, -2261, 7671, 3462, -7131, -4574, 6419, 5568, -5560, -6426, 4571, 7126, -3483, -7658, 2317, 8009, -1108, -8177, -123, 8157, 1341, -7959, -2525, 7583, 3645, -7047, -4682, 6360, 5611, -5544, -6417, 4613, 7083, -3594, -7600, 2505, 7957, -1373, -8153, 219, 8183, 931, -8053, -2058, 7765, 3137, -7332, -4150, 6759, 5078, -6065, -5906, 5261, 6619, -4367, -7208, 3398, 7663, -2376, -7980, 1317, 8153, -243, -8186, -830, 8077, 1880, -7834, -2894, 7460, 3852, -6968, -4742, 6364, 5548, -5664, -6262, 4878, 6871, -4022, -7372, 3109, 7755, -2156, -8020, 1176, 8162, -187, -8186, -800, 8089, 1767, -7879, -2703, 7559, 3594, -7137, -4430, 6620, 5199, -6019, -5894, 5340, 6505, -4599, -7029, 3802, 7457, -2964, -7790, 2094, 8022, -1206, -8156, 309, 8189, 583, -8127, -1464, 7968, 2318, -7721, -3142, 7387, 3922, -6975, -4654, 6488, 5328, -5938, -5942, 5326, 6486, -4666, -6960, 3962, 7358, -3226, -7681, 2462, 7924, -1682, -8090, 891, 8176, -100, -8186, -687, 8120, 1459, -7983, -2212, 7774, 2938, -7502, -3634, 7166, 4291, -6775, -4908, 6330, 5477, -5840, -5999, 5306, 6467, -4738, -6883, 4137, 7241, -3513, -7544, 2868, 7787, -2210, -7974, 1541, 8101, -870, -8174, 198, 8189, 466, -8153, -1123, 8062, 1763, -7924, -2387, 7736, 2989, -7505, -3568, 7231, 4118, -6920, -4640, 6572, 5129, -6193, -5586, 5783, 6006, -5349, -6392, 4891, 6739, -4416, -7050, 3922, 7321, -3418, -7557, 2902, 7753, -2381, -7913, 1854, 8034, -1328, -8122, 801, 8173, -279, -8191, -238, 8176, 746, -8130, -1247, 8054, 1733, -7950, -2209, 7818, 2669, -7663, -3114, 7483, 3541, -7283, -3953, 7061, 4344, -6823, -4718, 6566, 5070, -6296, -5404, 6011, 5717, -5717, -6011, 5410, 6283, -5097, -6537, 4775, 6769, -4448, -6983, 4116, 7175, -3782, -7351, 3445, 7507, -3108, -7646, 2770, 7766, -2435, -7871, 2100, 7959, -1770, -8033, 1442, 8090, -1120, -8135, 802, 8165, -491, -8185, 184, 8190, 114, -8187, -407, 8172, 690, -8149, -968, 8116, 1236, -8076, -1498, 8028, 1750, -7974, -1995, 7913, 2229, -7849, -2457, 7778, 2674, -7705, -2885, 7627, 3085, -7548, -3279, 7464, 3462, -7381, -3639, 7295, 3806, -7210, -3967, 7123, 4118, -7038, -4263, 6951, 4398, -6868, -4528, 6784, 4649, -6703, -4765, 6623, 4871, -6547, -4973, 6471, 5067, -6401, -5155, 6331, 5236, -6267, -5312, 6204, 5381, -6147, -5445, 6092, 5502, -6043, -5555, 5997, 5601, -5956, -5644, 5918, 5679, -5887, -5711, 5858, 5736, -5836, -5758, 5817, 5773, -5805, -5785, 5795, 5790, -5793, -5792, 5793, 5788, -5800, -5780, 5810, 5766, -5827, -5748, 5846, 5724, -5873, -5696, 5902, 5661, -5937, -5624, 5976, 5578, -6020, -5530, 6067, 5474, -6120, -5414, 6175, 5347, -6236, -5275, 6298, 5196, -6366, -5112, 6435, 5020, -6509, -4924, 6584, 4818, -6663, -4708, 6743, 4589, -6826, -4465, 6909, 4331, -6995, -4192, 7080, 4043, -7167, -3888, 7252, 3723, -7339, -3552, 7423, 3371, -7507, -3184, 7587, 2986, -7667, -2781, 7742, 2566, -7815, -2344, 7881, 2112, -7945, -1873, 8001, 1624, -8053, -1368, 8097, 1103, -8134, -831, 8161, 549, -8181, -261, 8190, -35, -8189, 337, 8176, -646, -8152, 960, 8114, -1281, -8063, 1605, 7997, -1936, -7917, 2267, 7820, -2603, -7709, 2939, 7578, -3277, -7432, 3613, 7265, -3950, -7082, 4283, 6877, -4613, -6655, 4936, 6412, -5255, -6150, 5565, 5866, -5866, -5563, 6155, 5239, -6434, -4896, 6696, 4532, -6945, -4151, 7174, 3748, -7386, -3330, 7576, 2893, -7745, -2441, 7887, 1972, -8006, -1492, 8095, 997, -8157, -493, 8187, -21, -8187, 540, 8151, -1065, -8083, 1591, 7978, -2119, -7838, 2643, 7659, -3162, -7444, 3672, 7190, -4172, -6899, 4656, 6569, -5124, -6204, 5569, 5799, -5992, -5362, 6386, 4888, -6751, -4383, 7080, 3845, -7374, -3282, 7626, 2690, -7836, -2078, 7999, 1444, -8114, -796, 8177, 134, -8189, 534, 8144, -1207, -8045, 1876, 7887, -2541, -7673, 3193, 7399, -3829, -7069, 4441, 6681, -5027, -6240, 5578, 5743, -6091, -5198, 6558, 4603, -6978, -3967, 7341, 3289, -7647, -2579, 7886, 1837, -8061, -1075, 8162, 293, -8191, 495, 8142, -1288, -8017, 2074, 7811, -2848, -7529, 3598, 7168, -4320, -6732, 5002, 6221, -5640, -5643, 6221, 4997, -6742, -4294, 7191, 3536, -7565, -2735, 7856, 1893, -8060, -1025, 8170, 137, -8186, 758, 8101, -1653, -7919, 2532, 7635, -3389, -7255, 4206, 6778, -4978, -6210, 5688, 5555, -6330, -4823, 6890, 4018, -7361, -3155, 7732, 2238, -7999, -1286, 8151, 307, -8189, 682, 8105, -1669, -7903, 2637, 7577, -3573, -7136, 4458, 6579, -5282, -5917, 6026, 5154, -6680, -4306, 7229, 3379, -7664, -2393, 7972, 1358, -8149, -295, 8187, -782, -8085, 1850, 7838, -2894, -7453, 3891, 6929, -4826, -6277, 5676, 5504, -6428, -4625, 7062, 3651, -7567, -2604, 7928, 1498, -8138, -357, 8188, -799, -8075, 1944, 7798, -3058, -7361, 4114, 6767, -5092, -6030, 5967, 5159, -6722, -4175, 7335, 3093, -7793, -1939, 8080, 733, -8191, 494, 8115, -1718, -7856, 2908, 7413, -4039, -6796, 5080, 6014, -6008, -5087, 6795, 4030, -7424, -2871, 7873, 1633, -8131, -350, 8185, -950, -8035, 2232, 7676, -3464, -7120, 4612, 6373, -5646, -5456, 6534, 4388, -7253, -3197, 7779, 1912, -8096, -570, 8190, -797, -8057, 2146, 7696, -3443, -7115, 4647, 6325, -5724, -5350, 6637, 4212, -7362, -2945, 7869, 1582, -8144, -167, 8172, -1263, -7952, 2658, 7483, -3979, -6780, 5180, 5859, -6224, -4748, 7073, 3479, -7699, -2092, 8076, 629, -8191, 860, 8033, -2329, -7607, 3724, 6921, -5001, -5997, 6111, 4861, -7017, -3554, 7680, 2114, -8078, -594, 8189, -955, -8009, 2474, 7537, -3913, -6790, 5212, 5788, -6327, -4569, 7208, 3172, -7825, -1651, 8145, 59, -8158, 1541, 7854, -3089, -7245, 4521, 6347, -5783, -5196, 6819, 3831, -7588, -2309, 8051, 684, -8190, 973, 7992, -2599, -7463, 4121, 6619, -5479, -5494, 6609, 4130, -7463, -2585, 7998, 921, -8191, 788, 8025, -2472, -7507, 4050, 6651, -5457, -5497, 6622, 4088, -7493, -2490, 8025, 770, -8191, 990, 7976, -2714, -7390, 4314, 6452, -5719, -5206, 6855, 3704, -7668, -2021, 8112, 231, -8164, 1575, 7813, -3312, -7076, 4890, 5982, -6230, -4586, 7259, 2950, -7926, -1160, 8187, -698, -8030, 2525, 7452, -4229, -6485, 5715, 5171, -6906, -3580, 7732, 1789, -8147, 102, 8122, -1997, -7657, 3787, 6768, -5377, -5504, 6673, 3928, -7602, -2128, 8106, 200, -8155, 1744, 7736, -3597, -6875, 5248, 5610, -6601, -4017, 7572, 2181, -8102, -212, 8152, -1778, -7719, 3667, 6818, -5343, -5504, 6699, 3848, -7652, -1954, 8135, -70, -8119, 2094, 7594, -3996, -6593, 5651, 5170, -6954, -3416, 7817, 1436, -8182, 642, 8017, -2686, -7332, 4560, 6163, -6142, -4585, 7321, 2696, -8019, -623, 8179, -1500, -7790, 3527, 6868, -5322, -5477, 6756, 3703, -7730, -1669, 8169, -490, -8040, 2619, 7344, -4572, -6128, 6204, 4470, -7401, -2488, 8067, 320, -8154, 1877, 7646, -3945, -6578, 5728, 5021, -7095, -3089, 7937, 918, -8189, 1325, 7824, -3478, -6867, 5371, 5382, -6860, -3482, 7825, 1306, -8190, 976, 7916, -3190, -7024, 5158, 5574, -6727, -3680, 7764, 1486, -8185, 832, 7947, -3092, -7068, 5105, 5610, -6710, -3690, 7766, 1459, -8187, 897, 7926, -3187, -7006, 5215, 5492, -6811, -3512, 7832, 1226, -8191, 1169, 7848, -3472, -6828, 5480, 5213, -7019, -3140, 7946, 784, -8180, 1645, 7689, -3937, -6515, 5883, 4754, -7308, -2562, 8076, 131, -8117, 2317, 7415, -4561, -6034, 6391, 4091, -7636, -1766, 8174, -732, -7951, 3166, 6978, -5310, -5346, 6955, 3200, -7944, -744, 8173, -1791, -7618, 4158, 6322, -6130, -4410, 7507, 2059, -8153, 499, 7995, -3015, -7046, 5237, 5390, -6943, -3192, 7954, 665, -8166, 1934, 7548, -4344, -6161, 6315, 4136, -7643, -1681, 8182, -956, -7875, 3498, 6742, -5682, -4900, 7272, 2535, -8098, 103, 8063, -2738, -7168, 5085, 5499, -6892, -3234, 7955, 610, -8157, 2084, 7466, -4559, -5955, 6535, 3780, -7795, -1182, 8188, -1555, -7669, 4124, 6284, -6235, -4188, 7644, 1610, -8188, 1157, 7795, -3799, -6508, 6008, 4464, -7528, -1898, 8175, -896, -7869, 3590, 6636, -5870, -4619, 7459, 2047, -8166, 772, 7897, -3508, -6682, 5826, 4656, -7447, -2062, 8165, -790, -7890, 3550, 6644, -5882, -4579, 7491, 1940, -8176, 945, 7841, -3719, -6524, 6032, 4381, -7590, -1682, 8187, -1240, -7746, 4007, 6310, -6269, -4062, 7727, 1282, -8189, 1668, 7586, -4410, -5992, 6578, 3606, -7887, -742, 8156, -2229, -7344, 4908, 5549, -6939, -3008, 8041, 56, -8062, 2909, 6989, -5487, -4965, 7320, 2255, -8156, 768, 7870, -3693, -6497, 6112, 4217, -7687, -1345, 8188, -1723, -7543, 4553, 5831, -6747, -3291, 7986, 276, -8091, 2784, 7036, -5452, -4968, 7338, 2176, -8167, 936, 7808, -3920, -6310, 6334, 3882, -7824, -878, 8160, -2264, -7289, 5074, 5328, -7134, -2569, 8128, -584, -7902, 3654, 6479, -6178, -4071, 7765, 1036, -8171, 2162, 7323, -5036, -5346, 7136, 2536, -8136, 672, 7869, -3783, -6373, 6306, 3872, -7843, -757, 8143, -2486, -7153, 5339, 5019, -7346, -2081, 8178, -1200, -7697, 4292, 5969, -6697, -3271, 8015, 32, -8029, 3216, 6724, -5944, -4312, 7695, 1180, -8177, 2152, 7297, -5133, -5199, 7260, 2223, -8172, 1130, 7706, -4302, -5936, 6747, 3151, -8049, 176, 7975, -3480, -6533, 6190, 3959, -7838, -697, 8127, -2694, -7003, 5619, 4650, -7568, -1479, 8187, -1961, -7363, 5058, 5231, -7265, -2165, 8178, -1295, -7631, 4527, 5710, -6952, -2756, 8123, -704, -7824, 4040, 6097, -6647, -3254, 8039, -194, -7957, 3610, 6403, -6367, -3662, 7944, 232, -8045, 3245, 6639, -6122, -3985, 7851, 573, -8100, 2952, 6813, -5924, -4228, 7770, 828, -8133, 2734, 6932, -5778, -4394, 7710, 999, -8151, 2594, 7004, -5690, -4488, 7676, 1086, -8158, 2535, 7030, -5662, -4510, 7670, 1088, -8157, 2555, 7012, -5695, -4462, 7695, 1006, -8148, 2656, 6950, -5789, -4341, 7746, 840, -8127, 2837, 6841, -5939, -4147, 7821, 590, -8090, 3094, 6678, -6142, -3874, 7911, 254, -8028, 3425, 6456, -6390, -3520, 8007, -167, -7931, 3824, 6164, -6673, -3079, 8096, -673, -7785, 4284, 5794, -6979, -2548, 8164, -1259, -7577, 4796, 5334, -7292, -1921, 8190, -1921, -7290, 5345, 4775, -7593, -1199, 8156, -2651, -6905, 5913, 4106, -7859, -383, 8039, -3434, -6408, 6480, 3322, -8063, 522, 7813, -4254, -5780, 7018, 2418, -8178, 1503, 7455, -5086, -5010, 7496, 1397, -8170, 2544, 6940, -5899, -4087, 7877, 269, -8008, 3617, 6249, -6656, -3011, 8121, -949, -7659, 4687, 5367, -7313, -1789, 8187, -2227, -7095, 5710, 4287, -7820, -438, 8034, -3526, -6295, 6634, 3014, -8126, 1009, 7624, -4792, -5246, 7397, 1566, -8177, 2505, 6927, -5962, -3951, 7935, -19, -7926, 3988, 5925, -6962, -2430, 8181, -1687, -7333, 5380, 4619, -7711, -726, 8077, -3361, -6376, 6590, 3033, -8130, 1095, 7572, -4948, -5054, 7521, 1217, -8143, 2941, 6638, -6337, -3395, 8075, -748, -7692, 4697, 5276, -7412, -1462, 8163, -2749, -6746, 6231, 3523, -8055, 645, 7719, -4649, -5307, 7403, 1458, -8163, 2789, 6708, -6287, -3428, 8076, -793, -7662, 4802, 5145, -7500, -1212, 8134, -3063, -6524, 6495, 3102, -8131, 1185, 7503, -5150, -4782, 7679, 714, -8058, 3557, 6168, -6834, -2537, 8182, -1820, -7213, 5665, 4189, -7902, 33, 7883, -4253, -5606, 7256, 1712, -8176, 2679, 6734, -6303, -3342, 8102, -1029, -7547, 5104, 4788, -7694, -624, 8030, -3730, -6007, 6990, 2208, -8191, 2248, 6966, -6045, -3670, 8046, -726, -7650, 4909, 4961, -7628, -781, 8054, -3642, -6054, 6969, 2218, -8191, 2294, 6924, -6117, -3548, 8075, -920, -7567, 5110, 4733, -7736, -440, 7979, -3997, -5756, 7200, 1744, -8173, 2815, 6599, -6503, -2964, 8160, -1606, -7261, 5676, 4074, -7965, 401, 7737, -4757, -5059, 7606, 768, -8041, 3772, 5907, -7114, -1881, 8178, -2756, -6615, 6510, 2916, -8168, 1729, 7182, -5822, -3864, 8024, -719, -7615, 5070, 4712, -7769, -262, 7918, -4281, -5461, 7417, 1195, -8105, 3470, 6104, -6990, -2072, 8185, -2658, -6649, 6503, 2882, -8174, 1856, 7095, -5976, -3624, 8082, -1079, -7454, 5421, 4292, -7926, 334, 7729, -4853, -4890, 7715, 369, -7932, 4283, 5416, -7465, -1029, 8069, -3722, -5877, 7185, 1637, -8152, 3177, 6272, -6888, -2197, 8187, -2657, -6612, 6580, 2703, -8187, 2165, 6897, -6273, -3159, 8155, -1708, -7136, 5971, 3564, -8104, 1287, 7331, -5683, -3922, 8036, -907, -7492, 5412, 4232, -7962, 566, 7619, -5166, -4500, 7884, -269, -7722, 4944, 4724, -7809, 14, 7799, -4754, -4910, 7739, 197, -7860, 4593, 5056, -7680, -366, 7902, -4468, -5169, 7632, 490, -7933, 4376, 5244, -7599, -573, 7950, -4323, -5288, 7581, 611, -7958, 4303, 5297, -7580, -607, 7954, -4323, -5275, 7594, 559, -7942, 4377, 5217, -7625, -469, 7916, -4469, -5127, 7669, 334, -7879, 4594, 5001, -7728, -157, 7825, -4755, -4839, 7795, -64, -7755, 4946, 4637, -7870, 327, 7662, -5168, -4396, 7947, -634, -7546, 5414, 4111, -8023, 982, 7398, -5686, -3782, 8091, -1372, -7217, 5973, 3404, -8148, 1800, 6995, -6275, -2979, 8182, -2265, -6730, 6582, 2502) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L32C31_i
    );

    L32C32_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (134, 7798, 4876, -4668, -7873, -381, 7629, 5266, -4259, -7992, -851, 7448, 5606, -3872, -8076, -1275, 7264, 5898, -3513, -8133, -1654, 7083, 6147, -3186, -8167, -1987, 6910, 6357, -2893, -8185, -2275, 6750, 6530, -2636, -8191, -2519, 6607, 6671, -2418, -8190, -2720, 6485, 6782, -2240, -8185, -2878, 6386, 6866, -2102, -8178, -2995, 6312, 6924, -2006, -8172, -3072, 6265, 6959, -1951, -8169, -3108, 6245, 6970, -1938, -8168, -3104, 6254, 6959, -1968, -8171, -3060, 6290, 6924, -2039, -8177, -2976, 6353, 6866, -2151, -8183, -2851, 6442, 6783, -2305, -8189, -2684, 6555, 6672, -2499, -8191, -2475, 6689, 6531, -2732, -8187, -2223, 6843, 6358, -3004, -8172, -1926, 7011, 6149, -3310, -8141, -1585, 7189, 5900, -3651, -8090, -1197, 7373, 5608, -4021, -8012, -764, 7556, 5269, -4417, -7901, -285, 7731, 4879, -4834, -7750, 237, 7890, 4435, -5266, -7551, 802, 8025, 3934, -5705, -7298, 1405, 8125, 3374, -6143, -6984, 2043, 8182, 2753, -6570, -6600, 2709, 8184, 2072, -6975, -6142, 3394, 8119, 1332, -7345, -5604, 4089, 7978, 539, -7667, -4981, 4782, 7748, -304, -7925, -4273, 5459, 7420, -1185, -8103, -3478, 6104, 6984, -2095, -8187, -2600, 6698, 6434, -3018, -8160, -1645, 7221, 5764, -3936, -8007, -622, 7653, 4972, -4830, -7715, 453, 7971, 4062, -5673, -7272, 1563, 8154, 3039, -6441, -6670, 2684, 8181, 1916, -7105, -5907, 3790, 8032, 710, -7636, -4983, 4849, 7692, -555, -8003, -3908, 5826, 7151, -1849, -8180, -2696, 6683, 6402, -3135, -8140, -1371, 7382, 5450, -4373, -7864, 36, 7884, 4304, -5516, -7338, 1484, 8153, 2988, -6516, -6558, 2926, 8159, 1533, -7323, -5530, 4307, 7876, -18, -7888, -4271, 5567, 7293, -1611, -8168, -2814, 6644, 6407, -3182, -8127, -1204, 7477, 5233, -4661, -7742, 498, 8009, 3801, -5971, -7002, 2220, 8190, 2159, -7038, -5918, 3880, 7986, 374, -7788, -4518, 5387, 7378, -1472, -8160, -2853, 6649, 6370, -3282, -8106, -997, 7579, 4991, -4952, -7598, 956, 8100, 3296, -6372, -6637, 2895, 8152, 1368, -7439, -5253, 4698, 7702, -687, -8060, -3507, 6237, 6745, -2738, -8166, -1493, 7393, 5317, -4646, -7717, 663, 8059, 3489, -6264, -6712, 2813, 8157, 1372, -7454, -5192, 4796, 7645, -889, -8100, -3246, 6445, 6529, -3122, -8118, -1005, 7607, 4865, -5141, -7471, 1358, 8158, 2764, -6763, -6178, 3648, 8016, 386, -7822, -4319, 5653, 7155, -2067, -8191, -2034, 7174, 5618, -4370, -7799, 481, 8039, 3519, -6290, -6645, 2991, 8128, 1037, -7616, -4806, 5239, 7394, -1591, -8180, -2441, 6978, 5873, -4092, -7884, 223, 7993, 3692, -6186, -6719, 2903, 8136, 1066, -7617, -4777, 5293, 7349, -1723, -8187, -2248, 7097, 5684, -4349, -7787, 587, 8070, 3303, -6480, -6423, 3391, 8052, 473, -7826, -4225, 5802, 7000, -2457, -8175, -1445, 7486, 5010, -5102, -7438, 1567, 8181, 2313, -7087, -5669, 4404, 7751, -744, -8103, -3077, 6653, 6207, -3735, -7964, -3, 7962, 3733, -6215, -6642, 3110, 8094, 665, -7785, -4291, 5788, 6981, -2546, -8164, -1240, 7589, 4752, -5393, -7245, 2048, 8189, 1725, -7396, -5128, 5039, 7441, -1627, -8188, -2123, 7216, 5421, -4741, -7585, 1283, 8169, 2434, -7064, -5643, 4502, 7684, -1023, -8148, -2662, 6945, 5796, -4332, -7749, 844, 8128, 2807, -6869, -5889, 4230, 7782, -751, -8119, -2874, 6836, 5920, -4202, -7790, 740, 8118, 2860, -6852, -5894, 4245, 7769, -816, -8130, -2768, 6911, 5807, -4361, -7722, 973, 8148, 2593, -7016, -5659, 4545, 7641, -1217, -8171, -2338, 7155, 5443, -4796, -7522, 1540, 8187, 1996, -7327, -5156, 5106, 7352, -1946, -8189, -1569, 7516, 4788, -5469, -7126, 2425, 8160, 1052, -7713, -4334, 5871, 6827, -2976, -8089, -449, 7899, 3785, -6302, -6444, 3587, 7953, -244, -8057, -3137, 6741, 5960, -4249, -7737, 1018, 8161, 2382, -7170, -5365, 4940, 7415, -1867, -8190, -1523, 7559, 4645, -5644, -6972, 2772, 8112, 560, -7883, -3794, 6328, 6384, -3719, -7904, 493, 8105, 2807, -6964, -5638, 4675, 7533, -1624, -8191, -1689, 7509, 4718, -5608, -6978, 2800, 8102, 451, -7923, -3626, 6471, 6212, -3991, -7806, 879, 8155, 2363, -7218, -5229, 5144, 7266, -2270, -8164, -954, 7787, 4021, -6206, -6462, 3667, 7900, -572, -8125, -2607, 7106, 5380, -5010, -7332, 2157, 8170, 1013, -7778, -4027, 6219, 6430, -3737, -7873, 703, 8143, 2427, -7212, -5195, 5221, 7193, -2471, -8138, -634, 7896, 3640, -6512, -6115, 4191, 7703, -1275, -8187, -1819, 7500, 4646, -5751, -6810, 3192, 8008, -190, -8080, -2833, 7021, 5454, -4988, -7312, 2267, 8155, 759, -7874, -3676, 6514, 6083, -4269, -7658, 1448, 8190, 1560, -7619, -4355, 6023, 6557, -3628, -7883, 754, 8157, 2212, -7354, -4882, 5584, 6903, -3088, -8020, 194, 8089, 2718, -7113, -5273, 5221, 7144, -2665, -8097, -227, 8016, 3082, -6920, -5543, 4952, 7298, -2368, -8137, -508, 7957, 3312, -6792, -5702, 4788, 7381, -2202, -8154, -649, 7926, 3413, -6739, -5758, 4737, 7402, -2171, -8155, -650, 7930, 3385, -6764, -5715, 4799, 7362, -2275, -8143, -511, 7967, 3230, -6867, -5569, 4973, 7257, -2512, -8110, -233, 8030, 2943, -7039, -5314, 5252, 7077, -2879, -8043, 186, 8105, 2518, -7266, -4939, 5623, 6806, -3367, -7922, 744, 8168, 1950, -7526, -4429, 6069, 6421, -3964, -7721, 1437, 8190, 1234, -7789, -3770, 6562, 5900, -4650, -7407, 2254, 8135, 369, -8017, -2949, 7069, 5217, -5398, -6945, 3177, 7959, -641, -8164, -1956, 7543, 4348, -6167, -6299, 4176, 7616, -1778, -8176, -793, 7927, 3276, -6903, -5435, 5206, 7057, -3010, -7994, 527, 8157, 1997, -7540, -4327, 6205, 6237, -4288, -7555, 1970, 8158, 525, -7999, -2966, 7095, 5123, -5539, -6805, 3477, 7856, -1104, -8190, -1364, 7779, 3701, -6670, -5701, 4964, 7183, -2821, -8025, 433, 8153, 1985, -7566, -4225, 6317, 6088, -4524, -7420, 2344, 8107, 30, -8099, -2397, 7399, 4552, -6076, -6317, 4243, 7546, -2062, -8142, -287, 8059, 2603, -7313, -4700, 5967, 6405, -4140, -7586, 1980, 8148, 331, -8055, -2611, 7317, 4675, -6001, -6364, 4213, 7544, -2102, -8133, -169, 8085, 2419, -7414, -4477, 6173, 6184, -4466, -7417, 2422, 8083, -204, -8140, -2025, 7586, 4094, -6471, -5856, 4880, 7179, -2937, -7974, 783, 8184, 1418, -7804, -3513, 6862, 5348, -5435, -6798, 3625, 7761, -1567, -8177, -597, 8019, 2711, -7306, -4632, 6090, 6227, -4462, -7393, 2533, 8052, -441, -8168, -1676, 7734, 3672, -6788, -5421, 5394, 6804, -3652, -7739, 1675, 8165, 402, -8064, -2448, 7444, 4329, -6352, -5931, 4860, 7150, -3068, -7919, 1088, 8190, 950, -7955, -2926, 7229, 4713, -6067, -6210, 4538, 7324, -2742, -7996, 787, 8188, 1207, -7895, -3124, 7138, 4850, -5967, -6290, 4453, 7359, -2689, -8004, 775, 8188, 1174, -7910, -3052, 7187, 4750, -6066, -6181, 4612, 7263, -2911, -7945, 1054, 8190, 850, -7993, -2705, 7367, 4406, -6352, -5869, 5003, 7015, -3398, -7793, 1620, 8161, 234, -8109, -2071, 7640, 3793, -6787, -5320, 5593, 6571, -4126, -7492, 2457, 8038, -675, -8188, -1135, 7937, 2881, -7305, -4484, 6323, 5864, -5046, -6963, 3533, 7728, -1862, -8131, 109, 8154, 1641, -7804, -3310, 7097, 4821, -6073, -6110, 4778, 7119, -3278, -7810, 1637, 8153, 68, -8139, -1765, 7772, 3377, -7074, -4840, 6075, 6089, -4825, -7079, 3376, 7768, -1794, -8134, 143, 8162, 1505, -7859, -3088, 7238, 4537, -6332, -5802, 5176, 6830, -3823, -7587, 2324, 8044, -743, -8191, -861, 8022, 2424, -7552, -3891, 6798, 5203, -5795, -6319, 4581, 7196, -3207, -7809, 1720, 8135, -180, -8170, -1362, 7913, 2847, -7380, -4228, 6591, 5454, -5580, -6488, 4379, 7295, -3038, -7854, 1599, 8145, -115, -8167, -1368, 7919, 2798, -7416, -4132, 6674, 5325, -5724, -6346, 4596, 7160, -3330, -7748, 1966, 8093, -549, -8190, -880, 8036, 2273, -7644, -3593, 7024, 4799, -6203, -5861, 5202, 6745, -4059, -7433, 2803, 7904, -1476, -8153, 112, 8171, 1246, -7965, -2565, 7541, 3806, -6917, -4940, 6109, 5935, -5145, -6770, 4049, 7422, -2856, -7882, 1594, 8135, -300, -8184, -997, 8026, 2260, -7672, -3463, 7130, 4573, -6421, -5569, 5559, 6425, -4572, -7127, 3482, 7657, -2319, -8009, 1107, 8176, 121, -8159, -1342, 7958, 2524, -7585, -3646, 7046, 4681, -6361, -5611, 5543, 6416, -4615, -7083, 3593, 7599, -2506, -7958, 1373, 8152, -220, -8184, -932, 8052, 2057, -7767, -3137, 7331, 4149, -6761, -5078, 6065, 5905, -5263, -6619, 4367, 7207, -3400, -7663, 2376, 7979, -1318, -8154, 242, 8185, 829, -8078, -1881, 7833, 2893, -7462, -3852, 6967, 4740, -6366, -5548, 5664, 6261, -4879, -6872, 4022, 7371, -3110, -7755, 2155, 8019, -1177, -8163, 186, 8185, 799, -8090, -1767, 7878, 2702, -7560, -3594, 7137, 4429, -6621, -5200, 6018, 5893, -5341, -6506, 4598, 7028, -3803, -7458, 2964, 7789, -2095, -8023, 1206, 8155, -310, -8190, -584, 8126, 1462, -7969, -2319, 7721, 3141, -7388, -3922, 6975, 4653, -6490, -5329, 5937, 5940, -5328, -6486, 4666, 6959, -3963, -7359, 3225, 7680, -2463, -7925, 1681, 8089, -892, -8177, 99, 8185, 686, -8121, -1459, 7982, 2211, -7775, -2939, 7501, 3632, -7167, -4291, 6774, 4906, -6331, -5478, 5839, 5998, -5307, -6468, 4737, 6882, -4138, -7242, 3512, 7543, -2869, -7788, 2209, 7973, -1542, -8102, 869, 8173, -200, -8190, -467, 8152, 1121, -8063, -1764, 7923, 2386, -7737, -2990, 7505, 3567, -7232, -4119, 6919, 4639, -6573, -5129, 6192, 5585, -5784, -6007, 5349, 6391, -4892, -6740, 4415, 7049, -3924, -7322, 3418, 7556, -2904, -7753, 2381, 7912, -1856, -8035, 1327, 8121, -802, -8174, 279, 8190, 237, -8177, -747, 8130, 1245, -8055, -1734, 7949, 2208, -7819, -2669, 7663, 3113, -7484, -3542, 7282, 3951, -7062, -4344, 6822, 4716, -6567, -5071, 6296, 5403, -6013, -5718, 5716, 6010, -5411, -6284, 5096, 6536, -4776, -6769, 4448, 6982, -4117, -7176, 3781, 7350, -3446, -7508, 3107, 7645, -2771, -7767, 2434, 7870, -2101, -7960, 1769, 8032, -1443, -8091, 1120, 8134, -803, -8166, 490, 8184, -185, -8191, -115, 8186, 406, -8173, -691, 8148, 967, -8117, -1237, 8075, 1497, -8029, -1750, 7973, 1993, -7914, -2230, 7848, 2456, -7779, -2675, 7704, 2884, -7628, -3086, 7547, 3278, -7465, -3463, 7380, 3638, -7296, -3807, 7209, 3966, -7124, -4119, 7037, 4262, -6952, -4399, 6867, 4527, -6785, -4650, 6702, 4764, -6624, -4872, 6546, 4972, -6472, -5067, 6400, 5154, -6332, -5237, 6266, 5311, -6205, -5382, 6146, 5444, -6093, -5503, 6042, 5554, -5998, -5602, 5955, 5643, -5919, -5680, 5886, 5710, -5859, -5737, 5835, 5757, -5818, -5774, 5804, 5784, -5796, -5791, 5792, 5791, -5794, -5789, 5799, 5779, -5811, -5767, 5826, 5747, -5847, -5725, 5872, 5695, -5903, -5662, 5936, 5623, -5977, -5579, 6019, 5529, -6068, -5475, 6119, 5413, -6176, -5348, 6235, 5274, -6299, -5197, 6365, 5111, -6436, -5021, 6508, 4923, -6585, -4819, 6662, 4707, -6744, -4590, 6825, 4464, -6910, -4332, 6994, 4191, -7081, -4044, 7166, 3887, -7253, -3724, 7338, 3551, -7424, -3372, 7506, 3183, -7588, -2987, 7666, 2780, -7742, -2567, 7814, 2343, -7882, -2113, 7944, 1872, -8002, -1625, 8052, 1368, -8098, -1104, 8133, 830, -8162, -550, 8180, 261, -8191, 34, 8188, -337, -8177, 645, 8151, -961, -8115, 1280, 8062, -1606, -7998, 1934, 7917, -2268, -7821, 2602, 7708, -2940, -7579, 3276, 7431, -3614, -7266, 3949, 7081, -4283, -6878, 4612, 6655, -4937, -6413, 5254, 6149, -5565, -5867, 5865, 5563, -6156, -5240, 6433, 4896, -6697, -4533, 6944, 4150, -7175, -3750, 7385, 3329, -7577, -2894, 7744, 2440, -7888, -1973, 8005, 1491, -8096, -998, 8156, 493, -8188, 19, 8186, -540, -8152, 1064, 8082, -1592, -7979, 2118, 7837, -2643, -7660, 3161, 7443, -3673, -7191, 4171, 6898, -4656, -6570, 5123, 6203, -5570, -5801, 5991, 5361, -6387, -4889, 6750, 4382, -7081, -3847, 7373, 3281, -7627, -2691, 7835, 2077, -8000, -1445, 8113, 795, -8178, -135, 8188, -535, -8145, 1205, 8044, -1877, -7888, 2540, 7672, -3193, -7400, 3828, 7069, -4442, -6682, 5026, 6239, -5578, -5745, 6090, 5197, -6559, -4605, 6977, 3966, -7342, -3290, 7645, 2578, -7887, -1838, 8060, 1074, -8163, -295, 8190, -496, -8143, 1287, 8016, -2074, -7813, 2846, 7529, -3598, -7169, 4319, 6731, -5003, -6223, 5639, 5642, -6222, -4999, 6740, 4294, -7192, -3538, 7564, 2734, -7857, -1895, 8059, 1025, -8171, -138, 8185, -759, -8102, 1652, 7918, -2533, -7636, 3387, 7254, -4207, -6779, 4977, 6210, -5689, -5557, 6329, 4823, -6891, -4020, 7360, 3154, -7733, -2240, 7998, 1286, -8152, -308, 8188, -682, -8107, 1668, 7902, -2637, -7578, 3571, 7135, -4459, -6580, 5281, 5916, -6027, -5156, 6679, 4305, -7229, -3381, 7663, 2392, -7973, -1359, 8148, 294, -8188, 781, 8084, -1851, -7839, 2893, 7452, -3892, -6930, 4825, 6277, -5677, -5505, 6427, 4625, -7063, -3653, 7566, 2604, -7929, -1499, 8137, 357, -8189, 797, 8075, -1944, -7799, 3056, 7360, -4114, -6768, 5091, 6030, -5968, -5161, 6721, 4175, -7336, -3095, 7792, 1938, -8081, -735, 8190, -494, -8116, 1717, 7856, -2909, -7414, 4038, 6796, -5081, -6016, 6007, 5086, -6796, -4031, 7423, 2870, -7873, -1635, 8130, 350, -8186, 949, 8034, -2232, -7678, 3463, 7119, -4612, -6374, 5644, 5456, -6534, -4389, 7252, 3197, -7780, -1914, 8095, 570, -8191, 795, 8057, -2146, -7697, 3442, 7115, -4647, -6327, 5722, 5350, -6638, -4213, 7360, 2944, -7870, -1584, 8143, 166, -8173, 1261, 7951, -2658, -7484, 3977, 6780, -5180, -5860, 6223, 4748, -7073, -3480, 7698, 2092, -8076, -631, 8190, -860, -8034, 2327, 7606, -3724, -6922, 5000, 5997, -6112, -4863, 7015, 3553, -7681, -2115, 8077, 594, -8190, 953, 8008, -2474, -7538, 3911, 6789, -5212, -5789, 6325, 4569, -7209, -3173, 7823, 1651, -8146, -60, 8157, -1541, -7855, 3087, 7244, -4522, -6348, 5782, 5196, -6820, -3833, 7586, 2309, -8052, -686, 8189, -973, -7993, 2597, 7462, -4122, -6620, 5478, 5494, -6609, -4131, 7462, 2585, -7999, -923, 8190, -789, -8026, 2470, 7506, -4051, -6653, 5455, 5497, -6622, -4090, 7492, 2490, -8025, -772, 8190, -991, -7977, 2712, 7389, -4315, -6453, 5718, 5205, -6856, -3706, 7667, 2021, -8113, -233, 8163, -1575, -7814, 3311, 7076, -4890, -5984, 6228, 4586, -7260, -2952, 7925, 1160, -8188, 696, 8029, -2525, -7454, 4227, 6485, -5715, -5173, 6904, 3579, -7732, -1791, 8146, -102, -8123, 1995, 7656, -3787, -6769, 5375, 5504, -6673, -3930, 7601, 2128, -8107, -202, 8154, -1744, -7738, 3596, 6874, -5248, -5612, 6600, 4017, -7572, -2183, 8101, 212, -8154, 1777, 7718, -3667, -6819, 5342, 5504, -6699, -3850, 7650, 1954, -8136, 68, 8118, -2094, -7595, 3994, 6593, -5651, -5172, 6953, 3416, -7817, -1438, 8181, -642, -8018, 2684, 7331, -4560, -6164, 6141, 4585, -7322, -2698, 8017, 623, -8180, 1498, 7789, -3527, -6870, 5320, 5477, -6756, -3705, 7729, 1669, -8170, 488, 8039, -2619, -7345, 4570, 6128, -6204, -4472, 7399, 2489, -8068, -322, 8153, -1877, -7647, 3943, 6578, -5728, -5023, 7094, 3089, -7937, -920, 8188, -1325, -7825, 3476, 6866, -5371, -5384, 6859, 3482, -7826, -1308, 8189, -976, -7917, 3188, 7023, -5158, -5576, 6725, 3680, -7764, -1488, 8184, -832, -7949, 3090, 7068, -5105, -5612, 6708, 3690, -7767, -1461, 8186, -897, -7928, 3185, 7005, -5215, -5494, 6809, 3512, -7833, -1228, 8190, -1169, -7849, 3470, 6828, -5480, -5214, 7017, 3140, -7947, -786, 8179, -1645, -7690, 3935, 6515, -5883, -4756, 7306, 2562, -8077, -133, 8116, -2317, -7417, 4559, 6034, -6391, -4093, 7635, 1766, -8175, 730, 7950, -3166, -6980, 5308, 5346, -6956, -3202, 7943, 744, -8174, 1789, 7618, -4158, -6324, 6128, 4410, -7508, -2061, 8152, -498, -7996, 3013, 7046, -5237, -5392, 6941, 3193, -7955, -668, 8165, -1933, -7550, 4342, 6161, -6315, -4138, 7641, 1681, -8183, 954, 7874, -3498, -6744, 5681, 4901, -7272, -2538, 8097, -102, -8064, 2736, 7168, -5085, -5501, 6890, 3234, -7956, -613, 8157, -2084, -7468, 4557, 5955, -6536, -3782, 7794, 1183, -8189, 1553, 7668, -4123, -6286, 6233, 4188, -7645, -1612, 8187, -1156, -7797, 3796, 6508, -6008, -4466, 7527, 1899, -8176, 894, 7868, -3590, -6638, 5868, 4619, -7459, -2050, 8165, -772, -7899, 3506, 6682, -5826, -4658, 7445, 2063, -8166, 788, 7889, -3550, -6646, 5880, 4579, -7492, -1942, 8175, -944, -7842, 3717, 6524, -6032, -4384, 7588, 1682, -8188, 1237, 7745, -4007, -6312, 6268, 4062, -7727, -1284, 8188, -1668, -7587, 4408, 5992, -6578, -3608, 7886, 742, -8157, 2227, 7343, -4908, -5551, 6937, 3009, -8041, -58, 8061, -2908, -6991, 5485, 4965, -7320, -2258, 8155, -767, -7871, 3691, 6497, -6112, -4219, 7685, 1346, -8189, 1720, 7543, -4552, -5833, 6745, 3292, -7987, -278, 8091, -2783, -7038, 5450, 4968, -7338, -2178, 8166, -935, -7810, 3917, 6310, -6334, -3884, 7823, 879, -8161, 2261, 7288, -5074, -5330, 7132, 2569, -8129, 582, 7901, -3653, -6481, 6176, 4072, -7766, -1039, 8171, -2161, -7324, 5033, 5346, -7136, -2539, 8135, -671, -7871, 3781, 6373, -6306, -3874, 7842, 757, -8144, 2484, 7153, -5338, -5022, 7344, 2081, -8179, 1198, 7697, -4292, -5971, 6695, 3271, -8016, -35, 8028, -3216, -6726, 5942, 4312, -7696, -1183, 8176, -2151, -7299, 5131, 5199, -7260, -2226, 8171, -1130, -7708, 4299, 5936, -6747, -3153, 8048, -175, -7976, 3478, 6533, -6190, -3962, 7836, 698, -8128, 2691, 7003, -5619, -4653, 7566, 1480, -8188, 1958, 7363, -5058, -5233, 7263, 2166, -8179, 1292, 7631, -4526, -5712, 6950, 2757, -8124, 701, 7823, -4040, -6099, 6645, 3254, -8040, 191, 7956, -3610, -6405, 6365, 3662, -7945, -235, 8044, -3245, -6641, 6120, 3985, -7851, -575, 8100, -2951, -6815, 5922, 4228, -7770, -831, 8132, -2733, -6934, 5776, 4395, -7710, -1002, 8150, -2594, -7006, 5688, 4488, -7676, -1088, 8157, -2534, -7032, 5660, 4511, -7671, -1091, 8156, -2555, -7014, 5693, 4462, -7695, -1009, 8147, -2656, -6952, 5786, 4342, -7747, -843, 8126, -2836, -6843, 5937, 4147, -7821, -592, 8089, -3093, -6680, 6140, 3875, -7912, -256, 8027, -3424, -6458, 6387, 3521, -8008, 165, 7930, -3823, -6166, 6671, 3080, -8097, 670, 7785, -4284, -5796, 6977, 2548, -8164, 1256, 7577, -4795, -5337, 7290, 1922, -8191, 1918, 7289, -5344, -4777, 7591, 1200, -8158, 2648, 6905, -5913, -4109, 7857, 384, -8040, 3432, 6408, -6480, -3325, 8062, -521, -7814, 4252, 5780, -7018, -2421, 8177, -1502, -7456, 5084, 5010, -7496, -1400, 8169, -2543, -6942, 5897, 4088, -7877, -272, 8007, -3616, -6252, 6654, 3012, -8122, 946, 7659, -4686, -5370, 7311, 1790, -8188, 2224, 7095, -5710, -4290, 7819, 439, -8036, 3523, 6295, -6634, -3017, 8125, -1008, -7626, 4789, 5246, -7397, -1569, 8176, -2504, -6929, 5960, 3951, -7935, 16, 7925, -3987, -5927, 6960, 2431, -8182, 1684, 7333, -5379, -4622, 7710, 727, -8078, 3358, 6376, -6590, -3036, 8129, -1094, -7573, 4945, 5054, -7521, -1220, 8142, -2940, -6640, 6335, 3395, -8076, 744, 7692, -4696, -5279, 7410, 1463, -8165, 2746, 6746, -6231, -3526, 8053, -644, -7720, 4646, 5308, -7403, -1462, 8162, -2788, -6710, 6285, 3429, -8076, 790, 7662, -4801, -5148, 7498, 1213, -8135, 3060, 6525, -6495, -3105, 8130, -1184, -7505, 5148, 4782, -7679, -718, 8057, -3557, -6171, 6832, 2538, -8183, 1817, 7213, -5664, -4192, 7901, -31, -7885, 4250, 5607, -7256, -1716, 8175, -2678, -6737, 6301, 3343, -8103, 1026, 7547, -5103, -4790, 7692, 625, -8032, 3727, 6008, -6990, -2211, 8190, -2247, -6968, 6042, 3671, -8047, 723, 7650, -4908, -4964, 7626, 782, -8056, 3639, 6055, -6969, -2221, 8190, -2293, -6927, 6114, 3549, -8076, 917, 7567, -5109, -4736, 7734, 441, -7980, 3994, 5757, -7199, -1747, 8172, -2813, -6602, 6501, 2965, -8161, 1603, 7261, -5676, -4077, 7963, -400, -7739, 4754, 5060, -7607, -771, 8040, -3771, -5909, 7112, 1882, -8179, 2753, 6616, -6509, -2919, 8167, -1728, -7184, 5819, 3865, -8025, 715, 7614, -5069, -4715, 7767, 264, -7919, 4278, 5461, -7417, -1198, 8104, -3469, -6107, 6988, 2073, -8186, 2655, 6649, -6503, -2885, 8173, -1855, -7097, 5974, 3625, -8082, 1076, 7454, -5420, -4295, 7924, -333, -7731, 4851, 4891, -7715, -373, 7931, -4282, -5419, 7463, 1030, -8070, 3719, 5877, -7185, -1640, 8151, -3175, -6275, 6885, 2198, -8188, 2654, 6612, -6579, -2706, 8186, -2163, -6899, 6270, 3161, -8156, 1705, 7136, -5970, -3567, 8103, -1285, -7333, 5681, 3924, -8037, 903, 7492, -5411, -4235, 7961, -565, -7621, 5163, 4501, -7884, 266, 7721, -4943, -4727, 7808, -12, -7801, 4751, 4911, -7739, -200, 7860, -4592, -5059, 7679, 368, -7904, 4465, 5170, -7632, -494, 7933, -4375, -5247, 7598, 574, -7952, 4319, 5289, -7581, -614, 7958, -4302, -5300, 7578, 609, -7956, 4320, 5276, -7594, -562, 7941, -4376, -5220, 7623, 470, -7917, 4466, 5128, -7669, -337, 7878, -4593, -5004, 7726, 159, -7827, 4752, 4840, -7795, 61, 7755, -4945, -4640, 7868, -325, -7664, 5165, 4398, -7947, 631, 7546, -5413, -4114, 8022, -980, -7400, 5683, 3784, -8092, 1369, 7218, -5972, -3408, 8146, -1798, -6998, 6273, 2981, -8183, 2262, 6730, -6582, -2505) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L32C32_i
    );

    L32C33_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-132, -7798, -4879, 4665, 7873, 382, -7629, -5269, 4256, 7991, 852, -7448, -5609, 3869, 8076, 1277, -7264, -5901, 3510, 8132, 1655, -7082, -6150, 3183, 8166, 1988, -6909, -6359, 2889, 8184, 2276, -6749, -6533, 2633, 8190, 2520, -6607, -6673, 2415, 8189, 2721, -6484, -6784, 2237, 8183, 2880, -6385, -6868, 2099, 8177, 2997, -6311, -6926, 2002, 8171, 3073, -6264, -6961, 1948, 8168, 3109, -6245, -6972, 1935, 8167, 3105, -6253, -6961, 1964, 8170, 3062, -6289, -6927, 2035, 8175, 2977, -6352, -6869, 2148, 8182, 2852, -6441, -6785, 2302, 8188, 2686, -6554, -6674, 2496, 8190, 2477, -6689, -6534, 2729, 8186, 2224, -6842, -6361, 3000, 8171, 1928, -7010, -6152, 3307, 8141, 1586, -7189, -5903, 3647, 8089, 1199, -7373, -5611, 4018, 8012, 765, -7556, -5272, 4414, 7900, 287, -7731, -4882, 4831, 7749, -236, -7890, -4438, 5263, 7551, -801, -8025, -3937, 5702, 7298, -1404, -8126, -3377, 6141, 6984, -2042, -8183, -2756, 6568, 6601, -2707, -8185, -2075, 6973, 6143, -3393, -8121, -1336, 7343, 5605, -4088, -7979, -542, 7665, 4982, -4781, -7750, 300, 7923, 4274, -5459, -7422, 1182, 8102, 3479, -6103, -6986, 2092, 8186, 2601, -6697, -6436, 3015, 8159, 1646, -7221, -5766, 3933, 8007, 624, -7653, -4975, 4827, 7715, -451, -7972, -4065, 5671, 7272, -1561, -8155, -3042, 6439, 6671, -2683, -8182, -1919, 7103, 5908, -3789, -8033, -713, 7634, 4984, -4848, -7694, 552, 8002, 3909, -5825, -7153, 1845, 8178, 2697, -6683, -6405, 3132, 8139, 1372, -7382, -5452, 4370, 7864, -35, -7884, -4307, 5514, 7338, -1483, -8154, -2991, 6514, 6559, -2925, -8160, -1536, 7321, 5531, -4306, -7878, 15, 7886, 4272, -5566, -7295, 1608, 8166, 2815, -6644, -6410, 3179, 8126, 1205, -7477, -5236, 4658, 7741, -497, -8009, -3804, 5969, 7003, -2219, -8191, -2162, 7036, 5918, -3879, -7988, -377, 7787, 4519, -5386, -7380, 1469, 8159, 2854, -6649, -6373, 3279, 8105, 998, -7580, -4994, 4949, 7598, -955, -8101, -3299, 6370, 6638, -2894, -8153, -1371, 7437, 5253, -4697, -7703, 683, 8059, 3507, -6237, -6747, 2735, 8165, 1494, -7393, -5319, 4643, 7717, -662, -8059, -3492, 6262, 6712, -2812, -8158, -1375, 7453, 5193, -4795, -7647, 886, 8099, 3247, -6445, -6531, 3119, 8117, 1006, -7608, -4868, 5139, 7471, -1357, -8159, -2767, 6761, 6178, -3647, -8017, -389, 7821, 4319, -5653, -7157, 2064, 8190, 2035, -7174, -5621, 4367, 7799, -480, -8039, -3521, 6288, 6645, -2990, -8130, -1040, 7614, 4807, -5239, -7396, 1588, 8179, 2442, -6978, -5875, 4089, 7883, -222, -7993, -3695, 6184, 6719, -2902, -8137, -1069, 7616, 4777, -5292, -7351, 1720, 8186, 2249, -7097, -5686, 4346, 7787, -586, -8071, -3305, 6478, 6423, -3390, -8053, -476, 7824, 4225, -5802, -7002, 2454, 8174, 1446, -7486, -5013, 5099, 7438, -1566, -8182, -2315, 7085, 5670, -4403, -7752, 742, 8102, 3077, -6653, -6210, 3733, 7963, 4, -7962, -3736, 6213, 6642, -3110, -8095, -668, 7783, 4292, -5787, -6983, 2543, 8163, 1241, -7589, -4755, 5390, 7245, -2047, -8190, -1728, 7394, 5128, -5039, -7443, 1624, 8186, 2124, -7216, -5423, 4739, 7585, -1282, -8170, -2437, 7062, 5644, -4502, -7686, 1020, 8147, 2663, -6945, -5799, 4330, 7749, -843, -8129, -2810, 6867, 5889, -4230, -7784, 748, 8117, 2875, -6836, -5922, 4199, 7789, -739, -8119, -2862, 6850, 5894, -4244, -7771, 813, 8129, 2768, -6911, -5809, 4358, 7722, -973, -8149, -2595, 7014, 5659, -4544, -7642, 1214, 8170, 2338, -7155, -5445, 4794, 7521, -1539, -8188, -1998, 7325, 5156, -5105, -7354, 1943, 8188, 1570, -7516, -4790, 5466, 7126, -2424, -8162, -1055, 7712, 4335, -5871, -6828, 2974, 8088, 449, -7899, -3788, 6300, 6444, -3587, -7954, 242, 8055, 3138, -6741, -5962, 4246, 7736, -1017, -8162, -2385, 7168, 5365, -4940, -7417, 1864, 8189, 1524, -7560, -4647, 5642, 6972, -2772, -8114, -563, 7882, 3795, -6328, -6386, 3717, 7904, -493, -8105, -2809, 6962, 5638, -4674, -7535, 1621, 8190, 1690, -7509, -4721, 5606, 6977, -2800, -8104, -454, 7921, 3626, -6471, -6214, 3989, 7805, -879, -8156, -2366, 7216, 5229, -5144, -7267, 2268, 8163, 954, -7788, -4024, 6204, 6462, -3667, -7902, 569, 8124, 2607, -7107, -5382, 5008, 7332, -2157, -8171, -1016, 7777, 4027, -6219, -6432, 3735, 7872, -703, -8144, -2429, 7211, 5195, -5221, -7195, 2469, 8137, 635, -7896, -3642, 6511, 6115, -4191, -7705, 1273, 8186, 1819, -7500, -4648, 5749, 6810, -3191, -8009, 188, 8079, 2834, -7021, -5456, 4986, 7312, -2267, -8156, -761, 7873, 3677, -6514, -6085, 4267, 7657, -1448, -8191, -1563, 7617, 4355, -6023, -6559, 3626, 7882, -753, -8158, -2215, 7352, 4882, -5584, -6905, 3086, 8019, -193, -8090, -2720, 7111, 5274, -5221, -7145, 2663, 8097, 228, -8017, -3085, 6918, 5543, -4952, -7300, 2365, 8136, 509, -7958, -3315, 6790, 5702, -4788, -7383, 2200, 8153, 649, -7927, -3415, 6737, 5758, -4737, -7404, 2169, 8154, 650, -7931, -3388, 6763, 5715, -4799, -7364, 2273, 8142, 512, -7968, -3232, 6866, 5569, -4973, -7259, 2510, 8109, 233, -8031, -2945, 7038, 5314, -5252, -7079, 2876, 8042, -186, -8105, -2520, 7265, 4939, -5623, -6807, 3364, 7921, -744, -8168, -1953, 7524, 4429, -6069, -6423, 3962, 7720, -1437, -8191, -1237, 7787, 3771, -6563, -5902, 4648, 7407, -2254, -8136, -371, 8016, 2949, -7069, -5219, 5396, 6945, -3177, -7960, 638, 8163, 1956, -7543, -4350, 6165, 6299, -4176, -7617, 1775, 8175, 793, -7928, -3278, 6901, 5435, -5206, -7058, 3008, 7993, -527, -8157, -2000, 7539, 4327, -6205, -6239, 4286, 7555, -1970, -8159, -527, 7997, 2966, -7095, -5125, 5537, 6805, -3477, -7858, 1102, 8189, 1365, -7780, -3703, 6668, 5700, -4964, -7185, 2819, 8024, -433, -8154, -1988, 7564, 4225, -6317, -6090, 4522, 7419, -2343, -8108, -33, 8098, 2397, -7400, -4554, 6075, 6317, -4243, -7547, 2060, 8141, 287, -8060, -2605, 7311, 4700, -5967, -6407, 4138, 7586, -1980, -8149, -334, 8054, 2611, -7317, -4677, 6000, 6363, -4214, -7546, 2100, 8132, 169, -8086, -2421, 7413, 4477, -6173, -6186, 4464, 7417, -2422, -8084, 202, 8139, 2025, -7586, -4096, 6469, 5855, -4880, -7180, 2935, 7973, -783, -8185, -1420, 7803, 3513, -6863, -5350, 5434, 6798, -3625, -7762, 1565, 8176, 597, -8019, -2713, 7305, 4632, -6090, -6229, 4460, 7393, -2533, -8053, 439, 8167, 1676, -7734, -3674, 6786, 5420, -5394, -6805, 3650, 7738, -1675, -8166, -404, 8063, 2448, -7444, -4331, 6351, 5930, -4860, -7152, 3066, 7919, -1088, -8191, -952, 7954, 2926, -7230, -4715, 6065, 6209, -4538, -7325, 2740, 7996, -787, -8189, -1209, 7894, 3124, -7138, -4852, 5966, 6289, -4453, -7360, 2687, 8003, -776, -8189, -1176, 7909, 3051, -7187, -4752, 6065, 6180, -4612, -7264, 2909, 7944, -1055, -8191, -852, 7992, 2705, -7367, -4407, 6350, 5868, -5003, -7017, 3396, 7792, -1620, -8162, -236, 8108, 2071, -7641, -3795, 6786, 5319, -5594, -6573, 4124, 7492, -2457, -8039, 673, 8187, 1135, -7938, -2883, 7304, 4484, -6324, -5866, 5044, 6963, -3533, -7730, 1860, 8131, -109, -8155, -1643, 7802, 3310, -7097, -4823, 6071, 6110, -4779, -7121, 3276, 7809, -1637, -8154, -70, 8138, 1764, -7773, -3378, 7072, 4839, -6075, -6091, 4823, 7079, -3376, -7769, 1792, 8133, -143, -8163, -1507, 7858, 3088, -7239, -4539, 6331, 5802, -5176, -6831, 3821, 7587, -2324, -8046, 742, 8190, 861, -8023, -2426, 7551, 3890, -6798, -5205, 5794, 6319, -4582, -7198, 3205, 7808, -1720, -8136, 178, 8169, 1362, -7914, -2849, 7379, 4227, -6592, -5455, 5578, 6488, -4380, -7296, 3037, 7853, -1599, -8146, 113, 8166, 1368, -7920, -2799, 7414, 4132, -6674, -5327, 5722, 6345, -4596, -7161, 3329, 7748, -1966, -8094, 547, 8189, 879, -8037, -2274, 7643, 3593, -7025, -4801, 6201, 5860, -5203, -6746, 4057, 7432, -2803, -7906, 1474, 8152, -112, -8172, -1248, 7964, 2565, -7541, -3808, 6915, 4940, -6109, -5936, 5143, 6769, -4050, -7424, 2855, 7881, -1595, -8136, 298, 8183, 996, -8027, -2261, 7671, 3462, -7131, -4574, 6419, 5568, -5560, -6426, 4571, 7126, -3483, -7658, 2317, 8009, -1108, -8177, -123, 8157, 1341, -7959, -2525, 7583, 3645, -7047, -4682, 6360, 5611, -5544, -6417, 4613, 7083, -3594, -7600, 2505, 7957, -1373, -8153, 219, 8183, 931, -8053, -2058, 7765, 3137, -7332, -4150, 6759, 5078, -6065, -5906, 5261, 6619, -4367, -7208, 3398, 7663, -2376, -7980, 1317, 8153, -243, -8186, -830, 8077, 1880, -7834, -2894, 7460, 3852, -6968, -4742, 6364, 5548, -5664, -6262, 4878, 6871, -4022, -7372, 3109, 7755, -2156, -8020, 1176, 8162, -187, -8186, -800, 8089, 1767, -7879, -2703, 7559, 3594, -7137, -4430, 6620, 5199, -6019, -5894, 5340, 6505, -4599, -7029, 3802, 7457, -2964, -7790, 2094, 8022, -1206, -8156, 309, 8189, 583, -8127, -1464, 7968, 2318, -7721, -3142, 7387, 3922, -6975, -4654, 6488, 5328, -5938, -5942, 5326, 6486, -4666, -6960, 3962, 7358, -3226, -7681, 2462, 7924, -1682, -8090, 891, 8176, -100, -8186, -687, 8120, 1459, -7983, -2212, 7774, 2938, -7502, -3634, 7166, 4291, -6775, -4908, 6330, 5477, -5840, -5999, 5306, 6467, -4738, -6883, 4137, 7241, -3513, -7544, 2868, 7787, -2210, -7974, 1541, 8101, -870, -8174, 198, 8189, 466, -8153, -1123, 8062, 1763, -7924, -2387, 7736, 2989, -7505, -3568, 7231, 4118, -6920, -4640, 6572, 5129, -6193, -5586, 5783, 6006, -5349, -6392, 4891, 6739, -4416, -7050, 3922, 7321, -3418, -7557, 2902, 7753, -2381, -7913, 1854, 8034, -1328, -8122, 801, 8173, -279, -8191, -238, 8176, 746, -8130, -1247, 8054, 1733, -7950, -2209, 7818, 2669, -7663, -3114, 7483, 3541, -7283, -3953, 7061, 4344, -6823, -4718, 6566, 5070, -6296, -5404, 6011, 5717, -5717, -6011, 5410, 6283, -5097, -6537, 4775, 6769, -4448, -6983, 4116, 7175, -3782, -7351, 3445, 7507, -3108, -7646, 2770, 7766, -2435, -7871, 2100, 7959, -1770, -8033, 1442, 8090, -1120, -8135, 802, 8165, -491, -8185, 184, 8190, 114, -8187, -407, 8172, 690, -8149, -968, 8116, 1236, -8076, -1498, 8028, 1750, -7974, -1995, 7913, 2229, -7849, -2457, 7778, 2674, -7705, -2885, 7627, 3085, -7548, -3279, 7464, 3462, -7381, -3639, 7295, 3806, -7210, -3967, 7123, 4118, -7038, -4263, 6951, 4398, -6868, -4528, 6784, 4649, -6703, -4765, 6623, 4871, -6547, -4973, 6471, 5067, -6401, -5155, 6331, 5236, -6267, -5312, 6204, 5381, -6147, -5445, 6092, 5502, -6043, -5555, 5997, 5601, -5956, -5644, 5918, 5679, -5887, -5711, 5858, 5736, -5836, -5758, 5817, 5773, -5805, -5785, 5795, 5790, -5793, -5792, 5793, 5788, -5800, -5780, 5810, 5766, -5827, -5748, 5846, 5724, -5873, -5696, 5902, 5661, -5937, -5624, 5976, 5578, -6020, -5530, 6067, 5474, -6120, -5414, 6175, 5347, -6236, -5275, 6298, 5196, -6366, -5112, 6435, 5020, -6509, -4924, 6584, 4818, -6663, -4708, 6743, 4589, -6826, -4465, 6909, 4331, -6995, -4192, 7080, 4043, -7167, -3888, 7252, 3723, -7339, -3552, 7423, 3371, -7507, -3184, 7587, 2986, -7667, -2781, 7742, 2566, -7815, -2344, 7881, 2112, -7945, -1873, 8001, 1624, -8053, -1368, 8097, 1103, -8134, -831, 8161, 549, -8181, -261, 8190, -35, -8189, 337, 8176, -646, -8152, 960, 8114, -1281, -8063, 1605, 7997, -1936, -7917, 2267, 7820, -2603, -7709, 2939, 7578, -3277, -7432, 3613, 7265, -3950, -7082, 4283, 6877, -4613, -6655, 4936, 6412, -5255, -6150, 5565, 5866, -5866, -5563, 6155, 5239, -6434, -4896, 6696, 4532, -6945, -4151, 7174, 3748, -7386, -3330, 7576, 2893, -7745, -2441, 7887, 1972, -8006, -1492, 8095, 997, -8157, -493, 8187, -21, -8187, 540, 8151, -1065, -8083, 1591, 7978, -2119, -7838, 2643, 7659, -3162, -7444, 3672, 7190, -4172, -6899, 4656, 6569, -5124, -6204, 5569, 5799, -5992, -5362, 6386, 4888, -6751, -4383, 7080, 3845, -7374, -3282, 7626, 2690, -7836, -2078, 7999, 1444, -8114, -796, 8177, 134, -8189, 534, 8144, -1207, -8045, 1876, 7887, -2541, -7673, 3193, 7399, -3829, -7069, 4441, 6681, -5027, -6240, 5578, 5743, -6091, -5198, 6558, 4603, -6978, -3967, 7341, 3289, -7647, -2579, 7886, 1837, -8061, -1075, 8162, 293, -8191, 495, 8142, -1288, -8017, 2074, 7811, -2848, -7529, 3598, 7168, -4320, -6732, 5002, 6221, -5640, -5643, 6221, 4997, -6742, -4294, 7191, 3536, -7565, -2735, 7856, 1893, -8060, -1025, 8170, 137, -8186, 758, 8101, -1653, -7919, 2532, 7635, -3389, -7255, 4206, 6778, -4978, -6210, 5688, 5555, -6330, -4823, 6890, 4018, -7361, -3155, 7732, 2238, -7999, -1286, 8151, 307, -8189, 682, 8105, -1669, -7903, 2637, 7577, -3573, -7136, 4458, 6579, -5282, -5917, 6026, 5154, -6680, -4306, 7229, 3379, -7664, -2393, 7972, 1358, -8149, -295, 8187, -782, -8085, 1850, 7838, -2894, -7453, 3891, 6929, -4826, -6277, 5676, 5504, -6428, -4625, 7062, 3651, -7567, -2604, 7928, 1498, -8138, -357, 8188, -799, -8075, 1944, 7798, -3058, -7361, 4114, 6767, -5092, -6030, 5967, 5159, -6722, -4175, 7335, 3093, -7793, -1939, 8080, 733, -8191, 494, 8115, -1718, -7856, 2908, 7413, -4039, -6796, 5080, 6014, -6008, -5087, 6795, 4030, -7424, -2871, 7873, 1633, -8131, -350, 8185, -950, -8035, 2232, 7676, -3464, -7120, 4612, 6373, -5646, -5456, 6534, 4388, -7253, -3197, 7779, 1912, -8096, -570, 8190, -797, -8057, 2146, 7696, -3443, -7115, 4647, 6325, -5724, -5350, 6637, 4212, -7362, -2945, 7869, 1582, -8144, -167, 8172, -1263, -7952, 2658, 7483, -3979, -6780, 5180, 5859, -6224, -4748, 7073, 3479, -7699, -2092, 8076, 629, -8191, 860, 8033, -2329, -7607, 3724, 6921, -5001, -5997, 6111, 4861, -7017, -3554, 7680, 2114, -8078, -594, 8189, -955, -8009, 2474, 7537, -3913, -6790, 5212, 5788, -6327, -4569, 7208, 3172, -7825, -1651, 8145, 59, -8158, 1541, 7854, -3089, -7245, 4521, 6347, -5783, -5196, 6819, 3831, -7588, -2309, 8051, 684, -8190, 973, 7992, -2599, -7463, 4121, 6619, -5479, -5494, 6609, 4130, -7463, -2585, 7998, 921, -8191, 788, 8025, -2472, -7507, 4050, 6651, -5457, -5497, 6622, 4088, -7493, -2490, 8025, 770, -8191, 990, 7976, -2714, -7390, 4314, 6452, -5719, -5206, 6855, 3704, -7668, -2021, 8112, 231, -8164, 1575, 7813, -3312, -7076, 4890, 5982, -6230, -4586, 7259, 2950, -7926, -1160, 8187, -698, -8030, 2525, 7452, -4229, -6485, 5715, 5171, -6906, -3580, 7732, 1789, -8147, 102, 8122, -1997, -7657, 3787, 6768, -5377, -5504, 6673, 3928, -7602, -2128, 8106, 200, -8155, 1744, 7736, -3597, -6875, 5248, 5610, -6601, -4017, 7572, 2181, -8102, -212, 8152, -1778, -7719, 3667, 6818, -5343, -5504, 6699, 3848, -7652, -1954, 8135, -70, -8119, 2094, 7594, -3996, -6593, 5651, 5170, -6954, -3416, 7817, 1436, -8182, 642, 8017, -2686, -7332, 4560, 6163, -6142, -4585, 7321, 2696, -8019, -623, 8179, -1500, -7790, 3527, 6868, -5322, -5477, 6756, 3703, -7730, -1669, 8169, -490, -8040, 2619, 7344, -4572, -6128, 6204, 4470, -7401, -2488, 8067, 320, -8154, 1877, 7646, -3945, -6578, 5728, 5021, -7095, -3089, 7937, 918, -8189, 1325, 7824, -3478, -6867, 5371, 5382, -6860, -3482, 7825, 1306, -8190, 976, 7916, -3190, -7024, 5158, 5574, -6727, -3680, 7764, 1486, -8185, 832, 7947, -3092, -7068, 5105, 5610, -6710, -3690, 7766, 1459, -8187, 897, 7926, -3187, -7006, 5215, 5492, -6811, -3512, 7832, 1226, -8191, 1169, 7848, -3472, -6828, 5480, 5213, -7019, -3140, 7946, 784, -8180, 1645, 7689, -3937, -6515, 5883, 4754, -7308, -2562, 8076, 131, -8117, 2317, 7415, -4561, -6034, 6391, 4091, -7636, -1766, 8174, -732, -7951, 3166, 6978, -5310, -5346, 6955, 3200, -7944, -744, 8173, -1791, -7618, 4158, 6322, -6130, -4410, 7507, 2059, -8153, 499, 7995, -3015, -7046, 5237, 5390, -6943, -3192, 7954, 665, -8166, 1934, 7548, -4344, -6161, 6315, 4136, -7643, -1681, 8182, -956, -7875, 3498, 6742, -5682, -4900, 7272, 2535, -8098, 103, 8063, -2738, -7168, 5085, 5499, -6892, -3234, 7955, 610, -8157, 2084, 7466, -4559, -5955, 6535, 3780, -7795, -1182, 8188, -1555, -7669, 4124, 6284, -6235, -4188, 7644, 1610, -8188, 1157, 7795, -3799, -6508, 6008, 4464, -7528, -1898, 8175, -896, -7869, 3590, 6636, -5870, -4619, 7459, 2047, -8166, 772, 7897, -3508, -6682, 5826, 4656, -7447, -2062, 8165, -790, -7890, 3550, 6644, -5882, -4579, 7491, 1940, -8176, 945, 7841, -3719, -6524, 6032, 4381, -7590, -1682, 8187, -1240, -7746, 4007, 6310, -6269, -4062, 7727, 1282, -8189, 1668, 7586, -4410, -5992, 6578, 3606, -7887, -742, 8156, -2229, -7344, 4908, 5549, -6939, -3008, 8041, 56, -8062, 2909, 6989, -5487, -4965, 7320, 2255, -8156, 768, 7870, -3693, -6497, 6112, 4217, -7687, -1345, 8188, -1723, -7543, 4553, 5831, -6747, -3291, 7986, 276, -8091, 2784, 7036, -5452, -4968, 7338, 2176, -8167, 936, 7808, -3920, -6310, 6334, 3882, -7824, -878, 8160, -2264, -7289, 5074, 5328, -7134, -2569, 8128, -584, -7902, 3654, 6479, -6178, -4071, 7765, 1036, -8171, 2162, 7323, -5036, -5346, 7136, 2536, -8136, 672, 7869, -3783, -6373, 6306, 3872, -7843, -757, 8143, -2486, -7153, 5339, 5019, -7346, -2081, 8178, -1200, -7697, 4292, 5969, -6697, -3271, 8015, 32, -8029, 3216, 6724, -5944, -4312, 7695, 1180, -8177, 2152, 7297, -5133, -5199, 7260, 2223, -8172, 1130, 7706, -4302, -5936, 6747, 3151, -8049, 176, 7975, -3480, -6533, 6190, 3959, -7838, -697, 8127, -2694, -7003, 5619, 4650, -7568, -1479, 8187, -1961, -7363, 5058, 5231, -7265, -2165, 8178, -1295, -7631, 4527, 5710, -6952, -2756, 8123, -704, -7824, 4040, 6097, -6647, -3254, 8039, -194, -7957, 3610, 6403, -6367, -3662, 7944, 232, -8045, 3245, 6639, -6122, -3985, 7851, 573, -8100, 2952, 6813, -5924, -4228, 7770, 828, -8133, 2734, 6932, -5778, -4394, 7710, 999, -8151, 2594, 7004, -5690, -4488, 7676, 1086, -8158, 2535, 7030, -5662, -4510, 7670, 1088, -8157, 2555, 7012, -5695, -4462, 7695, 1006, -8148, 2656, 6950, -5789, -4341, 7746, 840, -8127, 2837, 6841, -5939, -4147, 7821, 590, -8090, 3094, 6678, -6142, -3874, 7911, 254, -8028, 3425, 6456, -6390, -3520, 8007, -167, -7931, 3824, 6164, -6673, -3079, 8096, -673, -7785, 4284, 5794, -6979, -2548, 8164, -1259, -7577, 4796, 5334, -7292, -1921, 8190, -1921, -7290, 5345, 4775, -7593, -1199, 8156, -2651, -6905, 5913, 4106, -7859, -383, 8039, -3434, -6408, 6480, 3322, -8063, 522, 7813, -4254, -5780, 7018, 2418, -8178, 1503, 7455, -5086, -5010, 7496, 1397, -8170, 2544, 6940, -5899, -4087, 7877, 269, -8008, 3617, 6249, -6656, -3011, 8121, -949, -7659, 4687, 5367, -7313, -1789, 8187, -2227, -7095, 5710, 4287, -7820, -438, 8034, -3526, -6295, 6634, 3014, -8126, 1009, 7624, -4792, -5246, 7397, 1566, -8177, 2505, 6927, -5962, -3951, 7935, -19, -7926, 3988, 5925, -6962, -2430, 8181, -1687, -7333, 5380, 4619, -7711, -726, 8077, -3361, -6376, 6590, 3033, -8130, 1095, 7572, -4948, -5054, 7521, 1217, -8143, 2941, 6638, -6337, -3395, 8075, -748, -7692, 4697, 5276, -7412, -1462, 8163, -2749, -6746, 6231, 3523, -8055, 645, 7719, -4649, -5307, 7403, 1458, -8163, 2789, 6708, -6287, -3428, 8076, -793, -7662, 4802, 5145, -7500, -1212, 8134, -3063, -6524, 6495, 3102, -8131, 1185, 7503, -5150, -4782, 7679, 714, -8058, 3557, 6168, -6834, -2537, 8182, -1820, -7213, 5665, 4189, -7902, 33, 7883, -4253, -5606, 7256, 1712, -8176, 2679, 6734, -6303, -3342, 8102, -1029, -7547, 5104, 4788, -7694, -624, 8030, -3730, -6007, 6990, 2208, -8191, 2248, 6966, -6045, -3670, 8046, -726, -7650, 4909, 4961, -7628, -781, 8054, -3642, -6054, 6969, 2218, -8191, 2294, 6924, -6117, -3548, 8075, -920, -7567, 5110, 4733, -7736, -440, 7979, -3997, -5756, 7200, 1744, -8173, 2815, 6599, -6503, -2964, 8160, -1606, -7261, 5676, 4074, -7965, 401, 7737, -4757, -5059, 7606, 768, -8041, 3772, 5907, -7114, -1881, 8178, -2756, -6615, 6510, 2916, -8168, 1729, 7182, -5822, -3864, 8024, -719, -7615, 5070, 4712, -7769, -262, 7918, -4281, -5461, 7417, 1195, -8105, 3470, 6104, -6990, -2072, 8185, -2658, -6649, 6503, 2882, -8174, 1856, 7095, -5976, -3624, 8082, -1079, -7454, 5421, 4292, -7926, 334, 7729, -4853, -4890, 7715, 369, -7932, 4283, 5416, -7465, -1029, 8069, -3722, -5877, 7185, 1637, -8152, 3177, 6272, -6888, -2197, 8187, -2657, -6612, 6580, 2703, -8187, 2165, 6897, -6273, -3159, 8155, -1708, -7136, 5971, 3564, -8104, 1287, 7331, -5683, -3922, 8036, -907, -7492, 5412, 4232, -7962, 566, 7619, -5166, -4500, 7884, -269, -7722, 4944, 4724, -7809, 14, 7799, -4754, -4910, 7739, 197, -7860, 4593, 5056, -7680, -366, 7902, -4468, -5169, 7632, 490, -7933, 4376, 5244, -7599, -573, 7950, -4323, -5288, 7581, 611, -7958, 4303, 5297, -7580, -607, 7954, -4323, -5275, 7594, 559, -7942, 4377, 5217, -7625, -469, 7916, -4469, -5127, 7669, 334, -7879, 4594, 5001, -7728, -157, 7825, -4755, -4839, 7795, -64, -7755, 4946, 4637, -7870, 327, 7662, -5168, -4396, 7947, -634, -7546, 5414, 4111, -8023, 982, 7398, -5686, -3782, 8091, -1372, -7217, 5973, 3404, -8148, 1800, 6995, -6275, -2979, 8182, -2265, -6730, 6582, 2502) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L32C33_i
    );

    L40_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (134, 7798, 4877, -4667, -7874, -385, 7626, 5273, -4249, -7995, -868, 7440, 5624, -3847, -8082, -1313, 7244, 5932, -3463, -8140, -1721, 7044, 6202, -3102, -8174, -2091, 6847, 6435, -2767, -8190, -2423, 6655, 6635, -2459, -8190, -2718, 6473, 6804, -2181, -8181, -2977, 6305, 6947, -1933, -8164, -3201, 6152, 7065, -1718, -8144, -3390, 6018, 7161, -1535, -8123, -3547, 5905, 7236, -1386, -8103, -3670, 5814, 7293, -1271, -8086, -3762, 5746, 7334, -1189, -8073, -3823, 5701, 7358, -1142, -8066, -3853, 5682, 7366, -1129, -8065, -3852, 5688, 7360, -1151, -8070, -3820, 5718, 7338, -1206, -8081, -3758, 5773, 7301, -1296, -8096, -3665, 5852, 7246, -1420, -8115, -3540, 5953, 7173, -1578, -8136, -3382, 6076, 7081, -1768, -8157, -3191, 6218, 6966, -1992, -8176, -2965, 6378, 6828, -2247, -8188, -2705, 6553, 6662, -2532, -8191, -2408, 6740, 6467, -2847, -8181, -2074, 6935, 6239, -3189, -8154, -1702, 7134, 5976, -3556, -8105, -1293, 7332, 5673, -3945, -8029, -845, 7525, 5329, -4352, -7921, -361, 7706, 4940, -4772, -7774, 159, 7868, 4503, -5202, -7584, 713, 8006, 4018, -5633, -7345, 1299, 8110, 3481, -6060, -7051, 1911, 8174, 2894, -6475, -6697, 2545, 8189, 2255, -6869, -6278, 3194, 8146, 1568, -7232, -5791, 3851, 8037, 834, -7553, -5233, 4507, 7854, 58, -7821, -4601, 5150, 7588, -752, -8025, -3896, 5770, 7233, -1589, -8152, -3120, 6352, 6783, -2442, -8191, -2275, 6881, 6233, -3299, -8129, -1370, 7343, 5581, -4144, -7957, -413, 7720, 4828, -4962, -7663, 585, 7997, 3975, -5732, -7242, 1608, 8157, 3030, -6436, -6687, 2639, 8184, 2002, -7050, -5996, 3655, 8064, 904, -7554, -5172, 4634, 7786, -245, -7925, -4219, 5550, 7341, -1423, -8142, -3150, 6374, 6725, -2605, -8185, -1979, 7077, 5937, -3759, -8038, -729, 7631, 4984, -4854, -7689, 573, 8007, 3879, -5853, -7131, 1894, 8181, 2642, -6719, -6363, 3196, 8131, 1298, -7415, -5393, 4439, 7840, -118, -7906, -4236, 5575, 7301, -1564, -8161, -2917, 6561, 6513, -2993, -8153, -1470, 7349, 5486, -4353, -7864, 61, 7897, 4242, -5587, -7285, 1624, 8167, 2813, -6640, -6418, 3159, 8130, 1245, -7457, -5281, 4601, 7767, -407, -7988, -3903, 5883, 7072, -2075, -8190, -2330, 6937, 6057, -3687, -8036, -623, 7702, 4747, -5162, -7509, 1147, 8122, 3188, -6421, -6614, 2896, 8156, 1444, -7389, -5373, 4533, 7780, -405, -7996, -3833, 5965, 6991, -2268, -8191, -2061, 7102, 5808, -4040, -7939, -142, 7863, 4279, -5615, -7230, 1818, 8183, 2474, -6888, -6083, 3703, 8020, 489, -7765, -4544, 5393, 7357, -1560, -8170, -2694, 6769, 6212, -3542, -8052, -637, 7722, 4638, -5320, -7393, 1495, 8166, 2723, -6761, -6212, 3557, 8045, 585, -7745, -4569, 5396, 7341, -1628, -8177, -2565, 6863, 6078, -3753, -7999, -335, 7827, 4330, -5620, -7195, 1954, 8189, 2212, -7066, -5803, 4118, 7893, -116, -7953, -3913, 5972, 6933, -2468, -8181, -1663, 7342, 5364, -4640, -7701, 764, 8085, 3298, -6430, -6526, 3156, 8108, 905, -7656, -4736, 5288, 7377, -1606, -8179, -2474, 6946, 5932, -3995, -7920, 58, 7949, 3886, -6022, -6872, 2617, 8167, 1422, -7465, -5111, 4941, 7549, -1220, -8151, -2794, 6776, 6125, -3767, -7976, -148, 7903, 4021, -5935, -6927, 2546, 8171, 1444, -7467, -5087, 4986, 7516, -1328, -8163, -2641, 6880, 5981, -3979, -7911, 145, 7981, 3716, -6185, -6706, 2947, 8127, 972, -7660, -4661, 5416, 7266, -1925, -8191, -2007, 7229, 5470, -4610, -7678, 937, 8125, 2943, -6721, -6150, 3789, 7954, -4, -7957, -3779, 6162, 6704, -2983, -8119, -863, 7710, 4510, -5579, -7146, 2205, 8186, 1653, -7408, -5141, 4990, 7486, -1474, -8179, -2363, 7071, 5675, -4415, -7741, 796, 8112, 2990, -6719, -6122, 3867, 7922, -183, -8008, -3538, 6365, 6489, -3359, -8046, -366, 7876, 4005, -6027, -6788, 2896, 8122, 844, -7735, -4402, 5712, 7024, -2490, -8167, -1253, 7593, 4727, -5432, -7210, 2140, 8186, 1591, -7462, -4989, 5192, 7349, -1854, -8191, -1862, 7347, 5189, -4999, -7451, 1631, 8187, 2064, -7258, -5335, 4855, 7519, -1475, -8183, -2200, 7195, 5426, -4766, -7560, 1383, 8178, 2269, -7166, -5466, 4729, 7572, -1360, -8178, -2275, 7168, 5454, -4750, -7560, 1402, 8180, 2213, -7203, -5393, 4824, 7519, -1513, -8186, -2087, 7268, 5278, -4954, -7451, 1688, 8190, 1893, -7363, -5110, 5132, 7348, -1931, -8190, -1634, 7479, 4883, -5360, -7209, 2235, 8177, 1303, -7614, -4595, 5629, 7023, -2602, -8145, -906, 7755, 4238, -5936, -6787, 3025, 8083, 436, -7897, -3813, 6268, 6488, -3502, -7981, 102, 8024, 3310, -6619, -6121, 4022, 7825, -708, -8126, -2729, 6972, 5673, -4580, -7604, 1376, 8183, 2065, -7316, -5138, 5159, 7301, -2102, -8182, -1321, 7629, 4507, -5749, -6905, 2872, 8100, 496, -7895, -3776, 6327, 6399, -3677, -7922, 399, 8087, 2940, -6875, -5775, 4495, 7625, -1359, -8185, -2003, 7363, 5021, -5307, -7194, 2364, 8159, 967, -7766, -4134, 6081, 6609, -3394, -7989, 150, 8049, 3112, -6790, -5861, 4419, 7646, -1333, -8185, -1967, 7393, 4941, -5407, -7114, 2551, 8136, 708, -7854, -3851, 6314, 6372, -3772, -7877, 633, 8129, 2600, -7097, -5419, 4946, 7379, -2024, -8181, -1211, 7702, 4251, -6026, -6627, 3416, 7970, -284, -8083, -2889, 6950, 5611, -4754, -7471, 1834, 8187, 1359, -7658, -4343, 5968, 6662, -3381, -7975, 287, 8086, 2842, -6988, -5544, 4847, 7413, -1990, -8181, -1159, 7735, 4129, -6151, -6489, 3664, 7891, -647, -8139, -2462, 7199, 5205, -5218, -7192, 2484, 8134, 602, -7907, -3599, 6544, 6073, -4251, -7679, 1354, 8188, 1728, -7539, -4562, 5826, 6747, -3297, -7983, 309, 8098, 2715, -7086, -5358, 5090, 7251, -2394, -8142, -629, 7908, 3558, -6592, -5997, 4376, 7612, -1569, -8191, -1448, 7658, 4262, -6094, -6498, 3712, 7857, -838, -8164, -2144, 7381, 4834, -5622, -6881, 3120, 8014, -213, -8092, -2719, 7107, 5288, -5198, -7165, 2614, 8106, 302, -7998, -3176, 6858, 5634, -4841, -7367, 2206, 8155, 703, -7905, -3520, 6652, 5885, -4562, -7505, 1901, 8178, 992, -7828, -3758, 6501, 6049, -4372, -7588, 1703, 8186, 1168, -7778, -3893, 6415, 6135, -4273, -7627, 1614, 8188, 1233, -7761, -3929, 6397, 6145, -4271, -7623, 1636, 8187, 1187, -7779, -3866, 6449, 6081, -4363, -7578, 1766, 8182, 1030, -7831, -3703, 6568, 5939, -4549, -7486, 2006, 8166, 761, -7910, -3437, 6748, 5714, -4822, -7339, 2351, 8129, 378, -8003, -3062, 6977, 5396, -5175, -7124, 2798, 8056, -117, -8096, -2573, 7241, 4974, -5595, -6826, 3338, 7928, -724, -8167, -1966, 7520, 4436, -6065, -6425, 3960, 7720, -1437, -8191, -1235, 7788, 3770, -6563, -5903, 4646, 7409, -2248, -8137, -383, 8013, 2966, -7058, -5239, 5373, 6964, -3139, -7971, 586, 8158, 2020, -7514, -4417, 6107, 6360, -4086, -7658, 1656, 8182, 933, -7889, -3425, 6807, 5570, -5054, -7161, 2804, 8040, -284, -8130, -2260, 7423, 4577, -5997, -6446, 3990, 7686, -1605, -8184, -932, 7895, 3372, -6855, -5488, 5163, 7077, -2988, -7995, 534, 8158, 1963, -7559, -4273, 6254, 6179, -4374, -7511, 2091, 8145, 377, -8031, -2807, 7183, 4974, -5684, -6687, 3672, 7790, -1335, -8191, -1119, 7855, 3466, -6822, -5500, 5183, 7042, -3092, -7960, 731, 8176, 1687, -7679, -3954, 6513, 5871, -4787, -7278, 2651, 8054, -293, -8141, -2086, 7532, 4280, -6287, -6109, 4512, 7417, -2363, -8103, 20, 8108, 2318, -7441, -4460, 6159, 6227, -4374, -7481, 2233, 8118, 83, -8096, -2389, 7415, 4495, -6141, -6237, 4375, 7473, -2265, -8113, -21, 8106, 2299, -7462, -4392, 6231, 6134, -4518, -7396, 2456, 8079, -211, -8139, -2048, 7571, 4142, -6427, -5917, 4795, 7237, -2806, -8008, 608, 8174, 1629, -7730, -3740, 6709, 5567, -5196, -6979, 3302, 7874, -1171, -8191, -1041, 7910, 3171, -7058, -5068, 5697, 6594, -3933, -7647, 1891, 8150, 279, -8077, -2425, 7433, 4394, -6271, -6052, 4673, 7284, -2756, -8009, 652, 8180, 1490, -7791, -3527, 6870, 5316, -5487, -6744, 3735, 7711, -1740, -8162, -369, 8066, 2446, -7438, -4358, 6319, 5977, -4790, -7202, 2951, 7954, -927, -8191, -1153, 7898, 3152, -7101, -4947, 5853, 6420, -4239, -7486, 2360, 8077, -340, -8163, -1698, 7739, 3623, -6839, -5322, 5520, 6687, -3868, -7643, 1983, 8130, 15, -8128, -2009, 7635, 3875, -6690, -5507, 5348, 6807, -3696, -7704, 1830, 8146, 136, -8114, -2091, 7611, 3918, -6672, -5517, 5352, 6794, -3733, -7684, 1905, 8136, 23, -8131, -1947, 7671, 3755, -6788, -5351, 5531, 6647, -3976, -7578, 2206, 8091, -324, -8167, -1573, 7802, 3377, -7023, -4999, 5870, 6348, -4413, -7362, 2726, 7984, -903, -8191, -963, 7972, 2772, -7344, -4435, 6341, 5866, -5020, -6996, 3448, 7769, -1708, -8152, -113, 8126, 1922, -7700, -3632, 6894, 5157, -5755, -6428, 4338, 7382, -2718, -7979, 970, 8190, 817, -8013, -2562, 7456, 4178, -6552, -5596, 5342, 6747, -3891, -7585, 2263, 8069, -537, -8185, -1209, 7926, 2893, -7313, -4444, 6372, 5789, -5153, -6875, 3707, 7652, -2104, -8093, 413, 8179, 1289, -7912, -2932, 7303, 4442, -6387, -5760, 5201, 6828, -3801, -7607, 2244, 8065, -601, -8188, -1063, 7972, 2676, -7432, -4177, 6589, 5502, -5486, -6602, 4164, 7433, -2682, -7969, 1097, 8185, 524, -8083, -2120, 7664, 3627, -6953, -4992, 5975, 6159, -4774, -7089, 3395, 7747, -1896, -8115, 328, 8178, 1244, -7940, -2767, 7409, 4182, -6613, -5442, 5578, 6499, -4348, -7322, 2966, 7880, -1486, -8159, -44, 8151, 1564, -7860, -3027, 7297, 4378, -6488, -5577, 5460, 6581, -4252, -7361, 2905, 7891, -1467, -8159, -15, 8155, 1490, -7887, -2913, 7363, 4234, -6605, -5417, 5637, 6420, -4496, -7220, 3215, 7788, -1841, -8113, 414, 8185, 1020, -8008, -2418, 7586, 3736, -6938, -4938, 6084, 5987, -5054, -6857, 3878, 7519, -2594, -7963, 1238, 8172, 146, -8149, -1522, 7891, 2848, -7415, -4090, 6730, 5212, -5864, -6187, 4837, 6986, -3685, -7594, 2436, 7993, -1128, -8178, -207, 8144, 1528, -7897, -2806, 7444, 4004, -6801, -5096, 5985, 6051, -5022, -6850, 3934, 7472, -2754, -7908, 1509, 8144, -234, -8181, -1043, 8018, 2287, -7665, -3473, 7128, 4570, -6427, -5556, 5576, 6406, -4602, -7106, 3524, 7639, -2372, -7997, 1170, 8171, 52, -8165, -1268, 7975, 2450, -7614, -3574, 7087, 4614, -6412, -5552, 5601, 6367, -4678, -7045, 3659, 7572, -2571, -7942, 1433, 8146, -273, -8186, -888, 8059, 2025, -7775, -3118, 7337, 4143, -6761, -5084, 6054, 5921, -5237, -6644, 4324, 7236, -3335, -7692, 2288, 8001, -1205, -8165, 104, 8178, 991, -8047, -2065, 7771, 3096, -7363, -4069, 6826, 4964, -6177, -5772, 5423, 6477, -4585, -7070, 3672, 7542, -2705, -7889, 1697, 8104, -669, -8190, -366, 8143, 1388, -7970, -2385, 7672, 3337, -7260, -4235, 6737, 5062, -6118, -5811, 5408, 6468, -4625, -7028, 3777, 7481, -2882, -7826, 1948, 8057, -994, -8175, 30, 8178, 928, -8071, -1869, 7853, 2777, -7533, -3646, 7114, 4459, -6606, -5212, 6014, 5891, -5350, -6494, 4622, 7009, -3842, -7437, 3017, 7769, -2163, -8008, 1286, 8147, -401, -8191, -485, 8138, 1358, -7994, -2211, 7758, 3033, -7438, -3818, 7037, 4553, -6563, -5237, 6019, 5858, -5417, -6415, 4760, 6899, -4060, -7311, 3321, 7644, -2555, -7901, 1767, 8075, -969, -8172, 166, 8187, 632, -8127, -1421, 7989, 2188, -7780, -2933, 7500, 3643, -7156, -4318, 6750, 4948, -6290, -5533, 5777, 6065, -5221, -6544, 4624, 6963, -3995, -7324, 3337, 7621, -2658, -7858, 1962, 8030, -1259, -8141, 549, 8188, 158, -8176, -860, 8101, 1548, -7971, -2222, 7783, 2872, -7545, -3500, 7255, 4097, -6920, -4663, 6539, 5192, -6122, -5684, 5666, 6135, -5180, -6545, 4665, 6909, -4127, -7231, 3567, 7504, -2993, -7734, 2405, 7914, -1810, -8051, 1209, 8140, -608, -8186, 8, 8185, 585, -8144, -1171, 8059, 1744, -7937, -2305, 7774, 2847, -7577, -3372, 7344, 3874, -7081, -4356, 6786, 4810, -6466, -5241, 6118, 5643, -5750, -6018, 5359, 6363, -4952, -6679, 4528, 6964, -4092, -7220, 3643, 7444, -3187, -7640, 2722, 7803, -2254, -7939, 1782, 8043, -1311, -8121, 839, 8168, -371, -8190, -94, 8184, 551, -8154, -1003, 8098, 1444, -8021, -1878, 7919, 2299, -7799, -2710, 7656, 3107, -7497, -3492, 7318, 3861, -7125, -4218, 6915, 4557, -6693, -4883, 6457, 5191, -6211, -5485, 5953, 5761, -5688, -6023, 5413, 6267, -5133, -6496, 4845, 6707, -4555, -6905, 4258, 7085, -3961, -7251, 3660, 7401, -3359, -7537, 3056, 7658, -2755, -7767, 2453, 7860, -2155, -7942, 1857, 8010, -1564, -8068, 1272, 8112, -987, -8148, 703, 8171, -426, -8186, 152, 8190, 114, -8188, -377, 8175, 632, -8156, -882, 8129, 1125, -8096, -1363, 8056, 1592, -8012, -1817, 7961, 2032, -7907, -2243, 7848, 2446, -7786, -2643, 7719, 2831, -7652, -3015, 7580, 3189, -7508, -3359, 7433, 3521, -7358, -3677, 7281, 3825, -7205, -3969, 7126, 4104, -7050, -4235, 6973, 4358, -6898, -4477, 6822, 4588, -6749, -4695, 6676, 4794, -6606, -4890, 6537, 4979, -6471, -5064, 6406, 5142, -6345, -5217, 6285, 5285, -6230, -5351, 6175, 5409, -6126, -5465, 6078, 5515, -6035, -5562, 5994, 5602, -5958, -5640, 5923, 5673, -5894, -5702, 5867, 5726, -5846, -5748, 5827, 5764, -5813, -5778, 5801, 5785, -5795, -5791, 5792, 5791, -5794, -5789, 5797, 5781, -5807, -5772, 5819, 5756, -5836, -5738, 5856, 5714, -5881, -5689, 5908, 5657, -5940, -5622, 5975, 5582, -6014, -5539, 6056, 5490, -6102, -5438, 6150, 5380, -6203, -5319, 6257, 5252, -6315, -5181, 6375, 5103, -6439, -5023, 6503, 4935, -6572, -4844, 6640, 4745, -6713, -4642, 6785, 4532, -6860, -4419, 6935, 4297, -7012, -4171, 7088, 4037, -7166, -3898, 7242, 3751, -7320, -3600, 7395, 3440, -7471, -3276, 7544, 3102, -7617, -2924, 7685, 2737, -7754, -2546, 7817, 2345, -7878, -2139, 7934, 1925, -7988, -1706, 8034, 1478, -8077, -1245, 8113, 1004, -8144, -758, 8166, 504, -8183, -247, 8190, -19, -8190, 288, 8179, -564, -8161, 844, 8131, -1129, -8092, 1417, 8040, -1711, -7978, 2005, 7902, -2304, -7815, 2603, 7714, -2906, -7600, 3207, 7470, -3510, -7328, 3810, 7169, -4111, -6997, 4407, 6808, -4701, -6604, 4990, 6383, -5274, -6147, 5551, 5894, -5822, -5626, 6083, 5340, -6336, -5040, 6576, 4722, -6806, -4390, 7021, 4041, -7224, -3679, 7409, 3301, -7579, -2911, 7729, 2506, -7862, -2091, 7972, 1662, -8063, -1225, 8129, 777, -8173, -324, 8190, -139, -8183, 604, 8147, -1075, -8086, 1546, 7994, -2019, -7875, 2488, 7725, -2955, -7546, 3415, 7336, -3869, -7097, 4311, 6825, -4742, -6525, 5157, 6193, -5558, -5834, 5936, 5445, -6296, -5029, 6629, 4586, -6938, -4118, 7216, 3625, -7465, -3113, 7680, 2578, -7861, -2027, 8003, 1459, -8107, -880, 8170, 289, -8191, 307, 8168, -909, -8102, 1510, 7988, -2109, -7830, 2700, 7624, -3283, -7374, 3849, 7075, -4399, -6733, 4925, 6345, -5427, -5915, 5898, 5442, -6336, -4932, 6734, 4383, -7093, -3803, 7405, 3189, -7671, -2551, 7884, 1887, -8044, -1206, 8145, 510, -8190, 194, 8172, -904, -8094, 1611, 7952, -2312, -7748, 2999, 7480, -3669, -7151, 4313, 6760, -4928, -6312, 5504, 5805, -6040, -5248, 6526, 4638, -6961, -3986, 7335, 3292, -7649, -2565, 7893, 1807, -8067, -1029, 8166, 234, -8190, 567, 8133, -1370, -7998, 2163, 7782, -2941, -7488, 3694, 7114, -4415, -6666, 5094, 6144, -5726, -5555, 6298, 4902, -6809, -4192, 7247, 3430, -7609, -2627, 7886, 1787, -8078, -924, 8176, 42, -8182, 844, 8089, -1727, -7901, 2593, 7614, -3435, -7235, 4237, 6762, -4994, -6203, 5690, 5560, -6320, -4844, 6870, 4059, -7336, -3218, 7705, 2327, -7976, -1402, 8138, 450, -8191, 511, 8130, -1473, -7956, 2418, 7667, -3335, -7268, 4208, 6760, -5026, -6152, 5773, 5447, -6439, -4659, 7011, 3793, -7481, -2868, 7836, 1890, -8073, -880, 8182, -152, -8164, 1184, 8013, -2205, -7732, 3194, 7321, -4137, -6789, 5013, 6137, -5812, -5381, 6514, 4526, -7110, -3591, 7583, 2586, -7927, -1533, 8130, 445, -8191, 655, 8101, -1750, -7865, 2817, 7481, -3838, -6957, 4791, 6298, -5659, -5517, 6422, 4625, -7066, -3640, 7574, 2578, -7937, -1462, 8142, 309, -8187, 854, 8064, -2007, -7778, 3122, 7328, -4179, -6725, 5152, 5975, -6023, -5098, 6767, 4105, -7371, -3021, 7815, 1864, -8093, -663, 8190, -560, -8107, 1775, 7840, -2956, -7395, 4074, 6776, -5104, -6000, 6018, 5078, -6798, -4035, 7418, 2889, -7866, -1671, 8124, 406, -8188, 873, 8050, -2138, -7715, 3353, 7184, -4492, -6472, 5520, 5591, -6414, -4566, 7145, 3417, -7696, -2176, 8047, 871, -8189, 461, 8113, -1788, -7821, 3070, 7315, -4276, -6610, 5368, 5719, -6319, -4668, 7096, 3481, -7680, -2194, 8048, 837, -8190, 547, 8096, -1923, -7770, 3247, 7214, -4482, -6447, 5589, 5483, -6536, -4355, 7289, 3089, -7827, -1727, 8127, 304, -8181, 1131, 7981, -2538, -7534, 3869, 6847, -5086, -5943, 6144, 4845, -7012, -3589, 7655, 2210, -8055, -757, 8190, -729, -8059, 2194, 7658, -3593, -7002, 4876, 6105, -6000, -5000, 6922, 3719, -7612, -2307, 8040, 808, -8191, 723, 8055, -2236, -7635, 3672, 6941, -4985, -5998, 6122, 4834, -7043, -3492, 7709, 2015, -8096, -461, 8184, -1117, -7969, 2657, 7453, -4104, -6656, 5399, 5602, -6495, -4332, 7343, 2888, -7912, -1330, 8174, -288, -8118, 1898, 7739, -3440, -7054, 4848, 6083, -6068, -4865, 7046, 3445, -7742, -1881, 8121, 232, -8169, 1429, 7877, -3038, -7257, 4523, 6327, -5825, -5129, 6881, 3707, -7649, -2123, 8088, 441, -8181, 1264, 7916, -2921, -7305, 4453, 6367, -5795, -5146, 6881, 3689, -7663, -2064, 8101, 338, -8174, 1407, 7872, -3094, -7209, 4643, 6208, -5982, -4917, 7044, 3390, -7781, -1701, 8150, -77, -8134, 1854, 7727, -3550, -6948, 5077, 5828, -6364, -4423, 7341, 2794, -7963, -1025, 8190, -802, -8012, 2593, 7429, -4261, -6473, 5716, 5184, -6887, -3628, 7707, 1880, -8135, -31, 8141, -1826, -7724, 3592, 6900, -5176, -5712, 6489, 4216, -7463, -2493, 8038, 629, -8185, 1272, 7888, -3112, -7162, 4785, 6041, -6202, -4586, 7279, 2871, -7957, -993, 8190, -947, -7967, 2838, 7291, -4575, -6201, 6054, 4752, -7193, -3028, 7919, 1122, -8190, 852, 7983, -2783, -7310, 4555, 6203, -6064, -4727, 7216, 2964, -7941, -1021, 8190, -991, -7948, 2946, 7220, -4730, -6052, 6227, 4507, -7346, -2683, 8013, 685, -8184, 1359, 7843, -3325, -7010, 5085, 5729, -6529, -4083, 7559, 2170, -8110, -115, 8138, -1955, -7641, 3902, 6644, -5601, -5212, 6935, 3431, -7817, -1421, 8182, -691, -8005, 2760, 7289, -4650, -6083, 6230, 4460, -7394, -2531, 8054, 423, -8166, 1717, 7713, -3747, -6728, 5519, 5269, -6913, -3441, 7823, 1364, -8187, 812, 7969, -2938, -7186, 4858, 5884, -6436, -4158, 7552, 2125, -8125, 65, 8106, -2257, -7496, 4288, 6332, -6009, -4698, 7287, 2710, -8028, -517, 8168, -1723, -7696, 3836, 6640, -5665, -5079, 7066, 3125, -7932, -929, 8188, -1346, -7814, 3521, 6832, -5428, -5316, 6914, 3379, -7862, -1173, 8190, -1133, -7872, 3353, 6924, -5311, -5422, 6847, 3478, -7835, -1250, 8190, -1086, -7881, 3337, 6925, -5321, -5400, 6870, 3424, -7857, -1162, 8190, -1204, -7843, 3473, 6835, -5457, -5251, 6983, 3217, -7922, -907, 8185, -1488, -7751, 3758, 6646, -5712, -4967, 7173, 2851, -8016, -484, 8158, -1933, -7586, 4183, 6342, -6070, -4535, 7421, 2319, -8115, 108, 8081, -2532, -7322, 4731, 5898, -6508, -3937, 7695, 1611, -8183, 866, 7919, -3270, -6926, 5376, 5288, -6989, -3156, 7952, 723, -8174, 1781, 7626, -4124, -6359, 6081, 4484, -7465, -2179, 8137, -340, -8033, 2831, 7153, -5055, -5580, 6792, 3461, -7874, -1002, 8186, -1563, -7696, 3977, 6445, -6006, -4556, 7440, 2207, -8138, 365, 8021, -2908, -7100, 5161, 5458, -6899, -3261, 7937, 727, -8170, 1886, 7565, -4312, -6183, 6296, 4157, -7635, -1698, 8182, -945, -7877, 3492, 6745, -5680, -4903, 7271, 2537, -8098, 101, 8063, -2735, -7170, 5080, 5505, -6886, -3246, 7951, 630, -8159, 2058, 7479, -4529, -5983, 6507, 3827, -7777, -1247, 8190, -1478, -7699, 4042, 6349, -6163, -4290, 7597, 1745, -8183, 1000, 7846, -3638, -6622, 5868, 4642, -7436, -2130, 8155, -632, -7942, 3324, 6812, -5641, -4894, 7306, 2402, -8126, 373, 7998, -3111, -6933, 5487, 5049, -7222, -2566, 8104, -227, -8026, 2997, 6989, -5416, -5115, 7187, 2621, -8098, 192, 8030, -2989, -6989, 5426, 5092, -7207, -2572, 8107, -271, -8012, 3084, 6927, -5523, -4983, 7278, 2413, -8131, 461, 7967, -3284, -6803, 5697, 4779, -7397, -2147, 8160, -763, -7889, 3580, 6607, -5946, -4479, 7550, 1768, -8186, 1174, 7762, -3971, -6331, 6255, 4071, -7727, -1275, 8188, -1694, -7574, 4444, 5957, -6612, -3550, 7905, 665, -8149, 2313, 7301, -4987, -5474, 6994, 2904, -8063, 60, 8039, -3024, -6924, 5579, 4861, -7378, -2131, 8166, -898, -7834, 3808, 6417, -6197, -4109, 7727, 1224, -8186, 1835, 7498, -4644, -5758, 6803, 3202, -8007, -192, 8078, -2854, -7002, 5496, 4925, -7359, -2140, 8168, -958, -7806, 3921, 6314, -6325, -3906, 7812, 925, -8166, 2195, 7325, -5000, -5410, 7073, 2694, -8109, 422, 7945, -3483, -6603, 6030, 4274, -7682, -1303, 8185, -1869, -7461, 4764, 5609, -6946, -2908, 8077, -242, -7983, 3358, 6670, -5967, -4335, 7664, 1329, -8187, 1886, 7444, -4815, -5549, 7001, 2786, -8102, 414, 7937, -3556, -6529, 6142, 4091, -7768, -1005, 8166, -2247, -7272, 5145, 5217, -7230, -2328, 8160, -940, -7784, 4061, 6152, -6533, -3527, 7951, 323, -8082, 2936, 6896, -5723, -4583, 7576, 1513, -8190, 1809, 7454, -4839, -5487, 7071, 2606, -8134, 712, 7842, -3918, -6240, 6471, 3588, -7943, -330, 8077, -2991, -6848, 5809, 4453, -7646, -1299, 8181, -2083, -7320, 5112, 5201, -7269, -2185, 8175, -1214, -7671, 4406, 5834, -6840, -2981, 8083, -399, -7917, 3712, 6361, -6380, -3685, 7926, 353, -8075, 3045, 6791, -5909, -4299, 7723, 1034, -8161, 2419, 7135, -5444, -4826, 7492, 1642, -8191, 1843, 7405, -5000, -5273, 7249, 2175, -8180, 1324, 7611, -4587, -5645, 7008, 2634, -8141, 867, 7766, -4215, -5950, 6781, 3021, -8087, 476, 7880, -3890, -6194, 6576, 3338, -8027, 151, 7960, -3618, -6384, 6401, 3589, -7970, -106, 8014, -3404, -6524, 6263, 3775, -7921, -295, 8050, -3248, -6620, 6165, 3899, -7887, -417, 8069, -3154, -6674, 6110, 3963, -7869, -470, 8077, -3123, -6688, 6100, 3968, -7871, -456, 8073, -3154, -6663, 6135, 3913, -7891, -373, 8057, -3248, -6597, 6215, 3797, -7927, -223, 8026, -3403, -6489, 6336, 3620, -7977, -5, 7978, -3617, -6336, 6496, 3379, -8035, 281, 7906, -3889, -6131, 6689, 3072, -8095, 634, 7803, -4213, -5871, 6908, 2695, -8148, 1053, 7661, -4585, -5548, 7144, 2247, -8183, 1537, 7470, -4998, -5155, 7387, 1725, -8189, 2081, 7220, -5442, -4686, 7625, 1128, -8153, 2679, 6899, -5907, -4135, 7842, 457, -8058, 3324, 6495, -6378, -3496, 8022, -284, -7889, 4004, 5997, -6838, -2766, 8145, -1091, -7629, 4706, 5396, -7268, -1944, 8190, -1953, -7262, 5410, 4682, -7644, -1034, 8137, -2856, -6772, 6095, 3851, -7942, -43, 7961, -3782, -6145, 6735, 2902, -8134, 1016, 7642, -4705, -5371, 7299, 1840, -8190, 2124, 7159, -5597, -4445, 7753, 677, -8083, 3254, 6497, -6420, -3369, 8062, -568, -7786, 4372, 5645, -7136, -2151, 8189, -1866, -7274, 5437, 4601, -7700, -813, 8099, -3179, -6533, 6401, 3371, -8067, 616, 7761, -4459, -5553, 7210, 1976, -8191, 2091, 7150, -5648, -4341, 7808, 448, -8033, 3558, 6255, -6684, -2914, 8140, -1162, -7559, 4950, 5075, -7498, -1310, 8155, -2792, -6751, 6190, 3630, -8021, 415, 7810, -4362, -5606, 7196, 1962, -8191, 2188, 7080, -5781, -4145, 7886, 134, -7955, 3915, 5959, -6953, -2414, 8184, -1767, -7281, 5490, 4471, -7780, -486, 8027, -3634, -6163, 6798, 2667, -8171, 1537, 7377, -5340, -4625, 7725, 636, -8054, 3527, 6228, -6751, -2732, 8166, -1504, -7386, 5337, 4612, -7736, -588, 8041, -3601, -6165, 6815, 2607, -8177, 1664, 7305, -5487, -4434, 7808, 340, -7987, 3850, 5964, -6985, -2292, 8189, -2020, -7126, 5774, 4079, -7928, 106, 7870, -4268, -5613, 7238, 1778, -8181, 2560, 6821, -6183, -3537, 8062, -753, -7662, 4833, 5085, -7545, -1060, 8110, -3274, -6361, 6674, 2787, -8168, 1589, 7314, -5514, -4355, 7852, 133, -7924, 4131, 5698, -7202, -1817, 8180, -2600, -6777, 6261, 3389, -8096, 993, 7557, -5090, -4797, 7692, 618, -8029, 3746, 5989, -7007, -2174, 8190, -2294, -6940, 6081, 3616, -8059, 791, 7624, -4967, -4904, 7654, 703, -8041, 3712, 6000, -7012, -2143, 8190, -2370, -6884, 6165, 3481, -8088, 987, 7541, -5159, -4687, 7753, 389, -7969, 4030, 5731, -7214, -1722, 8170, -2825, -6599, 6499, 2975, -8159, 1577, 7277, -5643, -4124, 7948, -326, -7766, 4676, 5144, -7562, -901, 8066, -3633, -6024, 7020, 2071, -8188, 2542, 6753, -6353, -3168, 8140, -1434, -7330, 5580, 4170, -7943, 331, 7754, -4732, -5068, 7609, 742, -8032, 3828, 5851, -7162, -1770, 8170, -2894, -6518, 6616, 2734, -8181, 1946, 7065, -5995, -3629, 8075, -1007, -7498, 5313, 4442, -7869, 86, 7818, -4592, -5172, 7573, 799, -8036, 3842, 5813, -7206, -1644, 8156, -3083, -6369, 6776, 2435, -8191, 2323, 6839, -6303, -3172, 8148, -1577, -7229, 5793, 3847, -8040, 849, 7542, -5262, -4463, 7874, -151, -7786, 4717, 5016, -7663, -515, 7964, -4170, -5511, 7414, 1142, -8088, 3626, 5946, -7138, -1731, 8159, -3096, -6328, 6841, 2274, -8190, 2581, 6657, -6534, -2777, 8183, -2090, -6940, 6220, 3234, -8148, 1623, 7178, -5908, -3651, 8088, -1186, -7379, 5601, 4024, -8013, 778, 7544, -5307, -4359, 7924, -405, -7681, 5026, 4654, -7830, 64, 7789, -4765, -4914, 7731, 240, -7877, 4524, 5138, -7636, -512, 7945, -4308, -5331, 7544, 747, -7998, 4116, 5492, -7461, -948, 8037, -3954, -5626, 7386, 1113, -8068, 3818, 5730, -7326, -1245, 8087, -3714, -5811, 7278, 1341, -8102, 3637, 5864, -7246, -1404, 8109, -3594, -5894, 7229, 1431, -8113, 3580, 5899, -7229, -1426, 8111, -3599, -5881, 7244, 1385, -8105, 3647, 5837, -7277, -1312, 8091, -3728, -5770, 7322, 1202, -8073, 3836, 5676, -7384, -1060, 8045, -3977, -5556, 7456, 881, -8009, 4144, 5406, -7540, -669, 7959, -4339, -5229, 7631, 420, -7896, 4559, 5018, -7728, -138, 7813, -4803, -4775, 7824, -181, -7710, 5067, 4495, -7920, 532, 7581, -5351, -4179, 8008, -919, -7424, 5647, 3822, -8086, 1336, 7231, -5955, -3427, 8144, -1785, -7003, 6267, 2987, -8182, 2259, 6731, -6581, -2505) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L40_i
    );

    L40C31_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-131, -7798, -4880, 4663, 7873, 387, -7626, -5276, 4246, 7995, 870, -7439, -5627, 3843, 8081, 1315, -7243, -5936, 3459, 8139, 1723, -7044, -6205, 3098, 8173, 2093, -6846, -6438, 2763, 8189, 2425, -6654, -6637, 2455, 8189, 2720, -6472, -6807, 2176, 8180, 2979, -6304, -6950, 1929, 8163, 3203, -6151, -7067, 1714, 8143, 3392, -6017, -7163, 1531, 8121, 3548, -5904, -7239, 1382, 8101, 3672, -5812, -7296, 1267, 8084, 3764, -5744, -7336, 1185, 8072, 3824, -5700, -7360, 1138, 8065, 3854, -5681, -7369, 1125, 8064, 3854, -5687, -7362, 1147, 8069, 3822, -5717, -7341, 1202, 8079, 3760, -5772, -7303, 1292, 8095, 3667, -5851, -7249, 1416, 8114, 3542, -5952, -7176, 1574, 8135, 3384, -6075, -7083, 1764, 8156, 3193, -6217, -6969, 1988, 8174, 2967, -6377, -6830, 2243, 8187, 2707, -6552, -6665, 2529, 8190, 2410, -6739, -6470, 2843, 8181, 2076, -6934, -6242, 3186, 8154, 1704, -7133, -5979, 3553, 8105, 1295, -7332, -5677, 3941, 8029, 847, -7525, -5332, 4348, 7920, 363, -7706, -4943, 4769, 7774, -157, -7868, -4507, 5198, 7584, -711, -8006, -4021, 5630, 7345, -1297, -8111, -3485, 6057, 7051, -1909, -8175, -2898, 6472, 6698, -2543, -8190, -2259, 6866, 6279, -3192, -8148, -1571, 7229, 5792, -3850, -8039, -838, 7551, 5234, -4505, -7856, -62, 7819, 4602, -5149, -7590, 748, 8023, 3898, -5769, -7235, 1585, 8151, 3121, -6351, -6785, 2438, 8190, 2277, -6881, -6236, 3295, 8129, 1372, -7343, -5584, 4141, 7956, 414, -7720, -4831, 4958, 7664, -583, -7998, -3979, 5729, 7242, -1607, -8158, -3034, 6433, 6687, -2637, -8185, -2005, 7048, 5997, -3654, -8066, -908, 7552, 5173, -4633, -7788, 241, 7923, 4221, -5549, -7343, 1420, 8141, 3151, -6373, -6727, 2601, 8184, 1981, -7077, -5940, 3756, 8038, 731, -7631, -4988, 4851, 7689, -571, -8008, -3883, 5850, 7131, -1892, -8182, -2645, 6716, 6364, -3195, -8132, -1301, 7413, 5394, -4437, -7842, 114, 7905, 4237, -5574, -7303, 1560, 8160, 2918, -6560, -6516, 2990, 8152, 1471, -7349, -5489, 4349, 7864, -59, -7897, -4245, 5584, 7285, -1622, -8168, -2817, 6638, 6419, -3157, -8131, -1249, 7455, 5282, -4600, -7769, 403, 7986, 3904, -5882, -7075, 2072, 8189, 2332, -6937, -6059, 3683, 8035, 624, -7702, -4750, 5159, 7509, -1146, -8122, -3192, 6419, 6614, -2895, -8157, -1448, 7386, 5374, -4532, -7782, 402, 7995, 3835, -5964, -6993, 2264, 8190, 2062, -7102, -5811, 4037, 7938, 144, -7864, -4282, 5612, 7230, -1816, -8184, -2477, 6886, 6083, -3702, -8021, -492, 7763, 4546, -5392, -7359, 1556, 8169, 2695, -6768, -6215, 3538, 8052, 639, -7722, -4642, 5317, 7393, -1494, -8167, -2726, 6759, 6213, -3556, -8046, -589, 7743, 4570, -5395, -7343, 1625, 8176, 2566, -6862, -6081, 3750, 7998, 337, -7827, -4333, 5617, 7195, -1952, -8190, -2216, 7063, 5804, -4117, -7895, 113, 7951, 3914, -5971, -6935, 2465, 8180, 1664, -7342, -5367, 4637, 7701, -763, -8086, -3302, 6427, 6527, -3154, -8109, -908, 7654, 4737, -5287, -7379, 1602, 8178, 2475, -6946, -5935, 3992, 7920, -57, -7949, -3889, 6019, 6872, -2616, -8168, -1425, 7463, 5112, -4940, -7551, 1217, 8150, 2795, -6775, -6128, 3764, 7976, 150, -7903, -4024, 5932, 6927, -2545, -8172, -1448, 7465, 5088, -4985, -7518, 1325, 8162, 2643, -6879, -5984, 3976, 7911, -144, -7981, -3719, 6183, 6706, -2945, -8128, -975, 7658, 4662, -5415, -7268, 1922, 8190, 2008, -7228, -5473, 4607, 7678, -935, -8126, -2946, 6719, 6151, -3788, -7956, 1, 7956, 3780, -6161, -6706, 2980, 8118, 865, -7710, -4512, 5576, 7146, -2204, -8187, -1656, 7406, 5142, -4989, -7488, 1471, 8178, 2364, -7070, -5677, 4412, 7741, -795, -8113, -2993, 6717, 6123, -3865, -7923, 179, 8006, 3539, -6365, -6492, 3355, 8045, 367, -7877, -4009, 6025, 6788, -2895, -8124, -847, 7734, 4403, -5711, -7026, 2487, 8166, 1255, -7593, -4730, 5430, 7210, -2139, -8187, -1594, 7460, 4990, -5191, -7351, 1851, 8190, 1863, -7347, -5192, 4996, 7451, -1629, -8188, -2067, 7256, 5336, -4854, -7521, 1471, 8182, 2201, -7195, -5428, 4763, 7560, -1382, -8179, -2272, 7164, 5467, -4728, -7574, 1357, 8177, 2276, -7167, -5457, 4747, 7560, -1401, -8181, -2216, 7201, 5394, -4823, -7521, 1510, 8185, 2089, -7268, -5281, 4951, 7451, -1687, -8191, -1897, 7361, 5111, -5132, -7350, 1928, 8189, 1635, -7479, -4885, 5358, 7209, -2234, -8178, -1307, 7612, 4596, -5629, -7025, 2599, 8145, 907, -7756, -4241, 5933, 6787, -3024, -8084, -439, 7896, 3814, -6268, -6490, 3499, 7981, -101, -8025, -3313, 6617, 6121, -4021, -7827, 705, 8125, 2730, -6972, -5675, 4577, 7604, -1375, -8184, -2068, 7314, 5139, -5159, -7303, 2099, 8181, 1322, -7629, -4509, 5747, 6905, -2871, -8101, -500, 7893, 3777, -6327, -6401, 3674, 7922, -398, -8088, -2943, 6873, 5776, -4494, -7627, 1356, 8184, 2004, -7363, -5023, 5304, 7194, -2363, -8161, -970, 7764, 4135, -6081, -6611, 3392, 7989, -149, -8050, -3115, 6788, 5862, -4418, -7648, 1330, 8184, 1968, -7393, -4943, 5405, 7114, -2550, -8138, -711, 7852, 3852, -6313, -6375, 3769, 7877, -632, -8129, -2603, 7095, 5419, -4946, -7381, 2021, 8180, 1212, -7702, -4254, 6024, 6627, -3415, -7972, 281, 8082, 2890, -6950, -5613, 4752, 7471, -1833, -8188, -1362, 7657, 4343, -5968, -6664, 3378, 7975, -286, -8087, -2845, 6986, 5544, -4846, -7415, 1987, 8180, 1160, -7735, -4132, 6149, 6489, -3663, -7892, 644, 8138, 2462, -7200, -5208, 5216, 7191, -2483, -8136, -605, 7906, 3599, -6544, -6075, 4248, 7678, -1353, -8189, -1731, 7538, 4563, -5825, -6749, 3295, 7983, -309, -8099, -2717, 7084, 5358, -5090, -7253, 2392, 8141, 629, -7909, -3561, 6590, 5997, -4375, -7614, 1566, 8190, 1449, -7658, -4264, 6092, 6499, -3711, -7859, 835, 8163, 2145, -7382, -4837, 5619, 6881, -3119, -8015, 210, 8090, 2720, -7107, -5290, 5196, 7165, -2614, -8107, -305, 7997, 3176, -6858, -5636, 4838, 7367, -2205, -8156, -706, 7904, 3521, -6652, -5887, 4560, 7504, -1900, -8179, -995, 7826, 3758, -6501, -6051, 4369, 7588, -1702, -8187, -1171, 7776, 3894, -6415, -6137, 4271, 7626, -1614, -8189, -1236, 7759, 3929, -6397, -6147, 4268, 7623, -1635, -8188, -1190, 7778, 3867, -6449, -6083, 4361, 7578, -1766, -8183, -1033, 7830, 3704, -6568, -5941, 4546, 7486, -2005, -8167, -763, 7908, 3437, -6748, -5716, 4820, 7339, -2351, -8130, -381, 8002, 3063, -6977, -5398, 5173, 7124, -2797, -8057, 114, 8095, 2574, -7242, -4976, 5593, 6826, -3338, -7929, 721, 8166, 1966, -7520, -4438, 6063, 6425, -3960, -7722, 1435, 8190, 1236, -7788, -3772, 6561, 5903, -4646, -7410, 2245, 8136, 384, -8013, -2969, 7056, 5239, -5372, -6966, 3137, 7971, -585, -8159, -2023, 7513, 4417, -6107, -6362, 4084, 7658, -1656, -8183, -935, 7887, 3426, -6807, -5572, 5052, 7160, -2803, -8041, 282, 8129, 2261, -7423, -4579, 5995, 6446, -3990, -7687, 1602, 8184, 932, -7896, -3375, 6853, 5488, -5163, -7078, 2986, 7995, -533, -8159, -1966, 7558, 4274, -6254, -6181, 4372, 7510, -2091, -8146, -379, 8030, 2808, -7183, -4976, 5682, 6687, -3671, -7791, 1332, 8190, 1120, -7856, -3468, 6820, 5501, -5183, -7043, 3090, 7960, -731, -8177, -1689, 7677, 3954, -6513, -5873, 4785, 7278, -2650, -8056, 291, 8140, 2086, -7532, -4282, 6285, 6109, -4512, -7419, 2361, 8102, -20, -8109, -2320, 7440, 4460, -6159, -6229, 4372, 7480, -2233, -8119, -86, 8094, 2390, -7416, -4497, 6139, 6236, -4375, -7474, 2263, 8112, 22, -8107, -2301, 7460, 4392, -6231, -6136, 4516, 7396, -2456, -8080, 208, 8138, 2048, -7571, -4144, 6425, 5917, -4795, -7238, 2803, 8008, -607, -8175, -1631, 7729, 3740, -6710, -5569, 5194, 6979, -3301, -7875, 1169, 8190, 1041, -7910, -3173, 7056, 5068, -5697, -6596, 3931, 7646, -1891, -8151, -281, 8076, 2425, -7433, -4396, 6269, 6052, -4673, -7285, 2754, 8009, -651, -8180, -1493, 7789, 3527, -6870, -5318, 5485, 6743, -3735, -7713, 1737, 8161, 370, -8067, -2449, 7437, 4358, -6319, -5979, 4788, 7202, -2951, -7955, 925, 8190, 1153, -7898, -3154, 7100, 4947, -5853, -6422, 4237, 7486, -2360, -8078, 338, 8162, 1698, -7740, -3625, 6838, 5322, -5520, -6689, 3865, 7642, -1982, -8132, -18, 8127, 2009, -7636, -3877, 6688, 5507, -5348, -6809, 3694, 7704, -1830, -8147, -139, 8113, 2092, -7611, -3920, 6670, 5517, -5352, -6796, 3731, 7683, -1905, -8137, -26, 8130, 1947, -7671, -3757, 6786, 5351, -5531, -6649, 3974, 7577, -2206, -8092, 322, 8166, 1573, -7803, -3379, 7021, 4999, -5871, -6350, 4411, 7361, -2726, -7986, 901, 8190, 963, -7973, -2774, 7343, 4435, -6342, -5867, 5018, 6996, -3448, -7770, 1706, 8151, 114, -8127, -1924, 7699, 3632, -6894, -5159, 5754, 6428, -4338, -7383, 2716, 7978, -970, -8191, -819, 8012, 2562, -7456, -4180, 6550, 5596, -5343, -6749, 3889, 7584, -2262, -8070, 535, 8183, 1209, -7927, -2895, 7312, 4444, -6373, -5791, 5151, 6874, -3707, -7653, 2102, 8092, -413, -8180, -1291, 7910, 2932, -7304, -4444, 6385, 5760, -5201, -6829, 3799, 7607, -2244, -8066, 599, 8187, 1063, -7973, -2678, 7430, 4177, -6590, -5503, 5484, 6602, -4164, -7435, 2680, 7968, -1097, -8186, -526, 8082, 2120, -7665, -3629, 6951, 4992, -5975, -6160, 4773, 7089, -3396, -7749, 1894, 8114, -328, -8178, -1246, 7938, 2767, -7410, -4184, 6611, 5441, -5578, -6501, 4347, 7321, -2966, -7881, 1484, 8159, 44, -8151, -1566, 7859, 3027, -7298, -4380, 6487, 5577, -5460, -6583, 4251, 7361, -2905, -7892, 1465, 8158, 15, -8156, -1492, 7886, 2912, -7363, -4236, 6603, 5416, -5637, -6422, 4494, 7219, -3215, -7789, 1839, 8112, -414, -8186, -1021, 8006, 2418, -7586, -3738, 6937, 4938, -6084, -5989, 5053, 6856, -3878, -7521, 2592, 7962, -1239, -8173, -147, 8147, 1522, -7892, -2850, 7413, 4090, -6731, -5214, 5862, 6186, -4838, -6988, 3683, 7594, -2436, -7994, 1126, 8178, 207, -8145, -1530, 7896, 2806, -7444, -4006, 6800, 5096, -5985, -6052, 5020, 6850, -3934, -7474, 2752, 7907, -1509, -8145, 232, 8180, 1043, -8019, -2289, 7664, 3473, -7129, -4572, 6426, 5556, -5577, -6408, 4600, 7106, -3524, -7640, 2370, 7996, -1170, -8172, -53, 8164, 1268, -7976, -2451, 7613, 3574, -7088, -4616, 6411, 5552, -5602, -6368, 4676, 7045, -3659, -7573, 2569, 7941, -1433, -8147, 272, 8185, 888, -8060, -2027, 7774, 3118, -7338, -4144, 6759, 5084, -6055, -5923, 5236, 6643, -4324, -7237, 3333, 7691, -2288, -8003, 1203, 8164, -104, -8179, -993, 8046, 2065, -7772, -3097, 7361, 4068, -6827, -4966, 6175, 5772, -5424, -6478, 4583, 7070, -3672, -7543, 2703, 7888, -1698, -8105, 668, 8189, 366, -8144, -1390, 7969, 2384, -7673, -3339, 7259, 4235, -6738, -5064, 6116, 5810, -5409, -6469, 4624, 7027, -3778, -7482, 2880, 7826, -1948, -8058, 992, 8175, -30, -8179, -929, 8070, 1868, -7854, -2779, 7532, 3645, -7114, -4460, 6605, 5211, -6014, -5892, 5349, 6493, -4622, -7010, 3840, 7436, -3018, -7770, 2161, 8007, -1286, -8148, 400, 8190, 484, -8139, -1359, 7993, 2211, -7759, -3034, 7437, 3817, -7037, -4555, 6561, 5236, -6020, -5859, 5415, 6414, -4760, -6900, 4058, 7310, -3321, -7646, 2554, 7900, -1768, -8076, 968, 8171, -166, -8188, -634, 8126, 1420, -7990, -2190, 7779, 2932, -7501, -3645, 7155, 4318, -6751, -4950, 6289, 5533, -5778, -6066, 5220, 6543, -4625, -6964, 3994, 7323, -3337, -7623, 2657, 7858, -1963, -8032, 1257, 8141, -549, -8189, -160, 8175, 859, -8102, -1550, 7970, 2221, -7784, -2874, 7544, 3499, -7255, -4098, 6918, 4662, -6540, -5193, 6120, 5684, -5667, -6136, 5179, 6544, -4665, -6910, 4126, 7230, -3568, -7505, 2992, 7733, -2406, -7916, 1809, 8050, -1210, -8141, 607, 8185, -9, -8186, -586, 8143, 1171, -8060, -1746, 7936, 2304, -7775, -2848, 7576, 3371, -7345, -3876, 7080, 4355, -6787, -4812, 6465, 5240, -6119, -5644, 5749, 6017, -5360, -6364, 4951, 6678, -4529, -6965, 4091, 7220, -3643, -7445, 3185, 7639, -2722, -7804, 2253, 7938, -1783, -8044, 1310, 8120, -839, -8169, 370, 8189, 93, -8185, -552, 8153, 1002, -8099, -1446, 8020, 1877, -7920, -2300, 7798, 2710, -7657, -3108, 7496, 3491, -7319, -3863, 7124, 4217, -6916, -4558, 6692, 4882, -6458, -5193, 6210, 5485, -5954, -5763, 5687, 6022, -5414, -6268, 5132, 6495, -4846, -6709, 4554, 6904, -4259, -7086, 3960, 7250, -3660, -7402, 3358, 7537, -3057, -7659, 2754, 7766, -2454, -7861, 2154, 7941, -1858, -8011, 1563, 8067, -1273, -8113, 985, 8147, -704, -8172, 425, 8185, -153, -8191, -115, 8187, 376, -8176, -633, 8155, 882, -8130, -1126, 8095, 1362, -8057, -1593, 8011, 1816, -7962, -2034, 7906, 2243, -7848, -2447, 7785, 2642, -7720, -2832, 7651, 3014, -7581, -3190, 7507, 3358, -7434, -3522, 7357, 3676, -7282, -3826, 7204, 3968, -7127, -4105, 7049, 4234, -6974, -4359, 6897, 4476, -6823, -4589, 6748, 4694, -6677, -4795, 6605, 4889, -6538, -4980, 6470, 5063, -6407, -5143, 6344, 5216, -6286, -5287, 6229, 5350, -6176, -5410, 6125, 5464, -6079, -5516, 6034, 5561, -5995, -5603, 5957, 5639, -5924, -5674, 5893, 5701, -5868, -5727, 5845, 5747, -5828, -5765, 5812, 5777, -5802, -5786, 5794, 5790, -5793, -5792, 5793, 5788, -5798, -5782, 5806, 5771, -5820, -5757, 5835, 5737, -5857, -5715, 5880, 5687, -5909, -5657, 5940, 5621, -5976, -5583, 6013, 5538, -6057, -5491, 6101, 5437, -6151, -5381, 6202, 5318, -6258, -5253, 6314, 5180, -6376, -5104, 6438, 5022, -6504, -4936, 6571, 4842, -6641, -4746, 6712, 4641, -6786, -4533, 6859, 4417, -6936, -4298, 7011, 4170, -7089, -4038, 7165, 3897, -7243, -3752, 7319, 3599, -7396, -3441, 7470, 3275, -7545, -3103, 7616, 2923, -7687, -2738, 7753, 2544, -7818, -2346, 7877, 2138, -7935, -1926, 7987, 1705, -8035, -1479, 8076, 1244, -8114, -1005, 8143, 757, -8167, -505, 8182, 245, -8191, 18, 8189, -289, -8180, 564, 8160, -845, -8132, 1129, 8091, -1418, -8041, 1710, 7977, -2006, -7903, 2303, 7814, -2604, -7714, 2905, 7599, -3208, -7471, 3509, 7327, -3811, -7170, 4110, 6996, -4408, -6808, 4700, 6603, -4991, -6384, 5274, 6146, -5552, -5895, 5821, 5625, -6084, -5341, 6335, 5039, -6577, -4723, 6805, 4389, -7022, -4042, 7223, 3678, -7410, -3302, 7578, 2910, -7730, -2507, 7861, 2089, -7973, -1663, 8062, 1224, -8130, -778, 8172, 322, -8191, 138, 8182, -605, -8148, 1074, 8085, -1547, -7995, 2018, 7874, -2489, -7726, 2955, 7545, -3416, -7337, 3868, 7095, -4312, -6826, 4742, 6524, -5159, -6194, 5557, 5833, -5938, -5446, 6295, 5028, -6630, -4586, 6937, 4117, -7217, -3626, 7465, 3111, -7681, -2578, 7860, 2026, -8004, -1460, 8106, 879, -8171, -290, 8190, -309, -8169, 909, 8101, -1511, -7989, 2109, 7829, -2701, -7625, 3282, 7372, -3850, -7076, 4399, 6732, -4927, -6345, 5427, 5914, -5899, -5443, 6335, 4931, -6735, -4384, 7092, 3801, -7406, -3190, 7670, 2549, -7885, -1887, 8043, 1205, -8146, -510, 8189, -196, -8173, 904, 8093, -1612, -7953, 2312, 7747, -3001, -7481, 3669, 7150, -4314, -6761, 4927, 6311, -5506, -5806, 6040, 5246, -6528, -4639, 6960, 3985, -7337, -3292, 7648, 2563, -7894, -1807, 8067, 1027, -8167, -234, 8189, -569, -8134, 1369, 7997, -2164, -7783, 2941, 7487, -3695, -7115, 4415, 6665, -5095, -6145, 5725, 5554, -6300, -4902, 6808, 4191, -7248, -3431, 7608, 2626, -7888, -1788, 8077, 922, -8177, -42, 8181, -845, -8090, 1726, 7900, -2594, -7615, 3434, 7234, -4239, -6762, 4993, 6202, -5692, -5561, 6319, 4843, -6871, -4060, 7335, 3216, -7706, -2328, 7975, 1400, -8139, -450, 8190, -513, -8131, 1473, 7955, -2419, -7668, 3335, 7267, -4209, -6761, 5026, 6150, -5774, -5447, 6439, 4657, -7012, -3794, 7480, 2866, -7837, -1891, 8072, 878, -8183, 151, 8163, -1186, -8014, 2205, 7731, -3195, -7322, 4136, 6787, -5015, -6138, 5812, 5379, -6516, -4527, 7109, 3590, -7584, -2587, 7926, 1531, -8131, -445, 8190, -657, -8102, 1750, 7864, -2818, -7482, 3838, 6956, -4792, -6298, 5659, 5516, -6423, -4625, 7066, 3639, -7575, -2578, 7936, 1460, -8143, -309, 8186, -856, -8065, 2007, 7777, -3124, -7328, 4179, 6723, -5154, -5976, 6022, 5096, -6768, -4106, 7370, 3019, -7817, -1865, 8092, 661, -8191, 560, 8106, -1776, -7840, 2956, 7393, -4075, -6776, 5104, 5998, -6020, -5078, 6797, 4033, -7419, -2889, 7865, 1669, -8125, -406, 8187, -875, -8051, 2138, 7714, -3355, -7184, 4491, 6471, -5521, -5592, 6413, 4564, -7146, -3417, 7695, 2174, -8048, -871, 8188, -463, -8113, 1787, 7820, -3071, -7316, 4275, 6609, -5370, -5720, 6319, 4667, -7098, -3482, 7680, 2192, -8049, -837, 8189, -549, -8097, 1923, 7769, -3248, -7215, 4482, 6445, -5590, -5484, 6535, 4353, -7290, -3089, 7826, 1725, -8128, -304, 8180, -1132, -7982, 2538, 7533, -3871, -6847, 5086, 5941, -6146, -4845, 7012, 3587, -7657, -2211, 8054, 755, -8191, 729, 8058, -2196, -7659, 3593, 7000, -4877, -6105, 5999, 4999, -6923, -3719, 7611, 2305, -8041, -808, 8190, -725, -8056, 2235, 7634, -3674, -6942, 4985, 5997, -6124, -4834, 7043, 3490, -7710, -2015, 8096, 460, -8185, 1117, 7968, -2659, -7454, 4104, 6655, -5401, -5602, 6495, 4330, -7345, -2888, 7912, 1328, -8175, 288, 8116, -1900, -7740, 3440, 7053, -4850, -6083, 6068, 4863, -7047, -3445, 7741, 1879, -8122, -232, 8168, -1431, -7878, 3038, 7255, -4525, -6328, 5824, 5127, -6883, -3707, 7648, 2121, -8089, -441, 8180, -1266, -7917, 2921, 7303, -4455, -6368, 5795, 5144, -6882, -3689, 7663, 2062, -8102, -338, 8173, -1409, -7872, 3094, 7207, -4645, -6208, 5982, 4915, -7046, -3390, 7780, 1698, -8151, 77, 8133, -1856, -7727, 3550, 6946, -5079, -5828, 6363, 4421, -7343, -2794, 7962, 1023, -8191, 802, 8010, -2595, -7430, 4261, 6471, -5718, -5184, 6887, 3626, -7708, -1880, 8134, 29, -8141, 1827, 7723, -3594, -6901, 5176, 5711, -6491, -4216, 7462, 2491, -8039, -629, 8184, -1274, -7888, 3112, 7161, -4787, -6041, 6202, 4584, -7281, -2871, 7956, 991, -8191, 947, 7966, -2840, -7291, 4575, 6199, -6056, -4752, 7193, 3026, -7920, -1122, 8189, -854, -7984, 2783, 7309, -4557, -6203, 6064, 4725, -7217, -2964, 7941, 1019, -8191, 991, 7947, -2949, -7221, 4730, 6050, -6228, -4507, 7346, 2680, -8014, -684, 8183, -1362, -7844, 3326, 7008, -5087, -5729, 6529, 4081, -7561, -2170, 8109, 113, -8139, 1955, 7640, -3904, -6644, 5601, 5210, -6937, -3431, 7817, 1419, -8183, 691, 8003, -2762, -7289, 4651, 6081, -6232, -4460, 7393, 2529, -8055, -423, 8164, -1720, -7714, 3747, 6726, -5521, -5269, 6913, 3439, -7825, -1364, 8186, -815, -7970, 2939, 7184, -4860, -5884, 6436, 4156, -7553, -2125, 8124, -67, -8107, 2257, 7495, -4290, -6332, 6009, 4696, -7289, -2710, 8027, 514, -8169, 1723, 7695, -3838, -6640, 5665, 5077, -7068, -3125, 7931, 926, -8189, 1347, 7813, -3523, -6832, 5428, 5314, -6916, -3378, 7862, 1170, -8191, 1134, 7871, -3355, -6924, 5311, 5420, -6848, -3477, 7835, 1248, -8191, 1086, 7880, -3339, -6925, 5321, 5398, -6872, -3424, 7856, 1160, -8191, 1205, 7842, -3476, -6836, 5457, 5249, -6985, -3217, 7921, 905, -8186, 1488, 7749, -3761, -6647, 5712, 4965, -7175, -2851, 8015, 482, -8159, 1933, 7584, -4185, -6342, 6070, 4533, -7423, -2318, 8114, -110, -8082, 2532, 7321, -4733, -5898, 6508, 3935, -7696, -1610, 8182, -869, -7920, 3271, 6924, -5378, -5288, 6989, 3154, -7953, -723, 8173, -1783, -7627, 4125, 6357, -6083, -4484, 7465, 2177, -8139, 341, 8032, -2833, -7153, 5055, 5578, -6794, -3461, 7873, 999, -8187, 1564, 7695, -3980, -6445, 6006, 4553, -7442, -2206, 8137, -368, -8022, 2909, 7098, -5163, -5458, 6899, 3259, -7939, -726, 8169, -1888, -7566, 4312, 6181, -6298, -4157, 7635, 1695, -8183, 945, 7876, -3494, -6745, 5680, 4900, -7273, -2536, 8097, -104, -8064, 2736, 7169, -5083, -5505, 6886, 3243, -7953, -629, 8158, -2061, -7480, 4529, 5981, -6509, -3826, 7776, 1244, -8191, 1479, 7697, -4044, -6349, 6163, 4288, -7598, -1744, 8182, -1002, -7846, 3639, 6620, -5870, -4642, 7436, 2128, -8156, 632, 7941, -3327, -6812, 5641, 4891, -7308, -2401, 8126, -375, -7998, 3111, 6931, -5489, -5048, 7222, 2563, -8105, 228, 8025, -3000, -6990, 5416, 5113, -7189, -2620, 8097, -195, -8030, 2990, 6987, -5429, -5092, 7207, 2569, -8108, 272, 8011, -3087, -6927, 5523, 4980, -7280, -2412, 8130, -463, -7967, 3284, 6802, -5699, -4778, 7396, 2145, -8161, 764, 7887, -3583, -6607, 5946, 4476, -7552, -1767, 8185, -1177, -7762, 3972, 6329, -6257, -4070, 7727, 1273, -8189, 1695, 7572, -4446, -5957, 6612, 3547, -7906, -664, 8147, -2316, -7301, 4988, 5472, -6996, -2904, 8062, -63, -8040, 3025, 6922, -5581, -4861, 7378, 2129, -8168, 899, 7832, -3810, -6416, 6197, 4107, -7729, -1223, 8185, -1837, -7498, 4644, 5756, -6805, -3202, 8006, 189, -8078, 2854, 7000, -5498, -4924, 7359, 2138, -8169, 959, 7804, -3924, -6313, 6325, 3903, -7814, -924, 8165, -2198, -7325, 5000, 5408, -7075, -2693, 8108, -425, -7946, 3484, 6601, -6032, -4273, 7682, 1300, -8186, 1870, 7460, -4767, -5609, 6946, 2905, -8078, 243, 7982, -3360, -6670, 5968, 4332, -7666, -1328, 8186, -1889, -7444, 4816, 5546, -7003, -2785, 8101, -417, -7937, 3556, 6527, -6145, -4090, 7767, 1002, -8167, 2248, 7270, -5148, -5216, 7230, 2325, -8161, 941, 7782, -4064, -6152, 6534, 3524, -7953, -322, 8081, -2938, -6896, 5723, 4580, -7578, -1512, 8189, -1812, -7454, 4840, 5485, -7073, -2605, 8133, -715, -7842, 3919, 6238, -6473, -3587, 7943, 327, -8078, 2992, 6845, -5811, -4452, 7645, 1296, -8182, 2084, 7318, -5115, -5200, 7269, 2182, -8177, 1215, 7670, -4409, -5834, 6840, 2978, -8085, 400, 7916, -3715, -6361, 6380, 3682, -7927, -352, 8074, -3048, -6791, 5909, 4296, -7724, -1033, 8160, -2422, -7135, 5445, 4824, -7494, -1641, 8190, -1846, -7405, 5000, 5270, -7251, -2174, 8179, -1327, -7612, 4588, 5643, -7010, -2633, 8141, -871, -7767, 4215, 5948, -6783, -3020, 8086, -479, -7880, 3891, 6192, -6578, -3337, 8026, -154, -7960, 3619, 6382, -6403, -3588, 7969, 103, -8015, 3405, 6522, -6265, -3774, 7921, 292, -8050, 3249, 6618, -6167, -3898, 7886, 413, -8070, 3155, 6672, -6112, -3962, 7869, 467, -8077, 3124, 6686, -6103, -3967, 7870, 452, -8073, 3155, 6660, -6138, -3912, 7890, 370, -8057, 3249, 6595, -6218, -3796, 7927, 220, -8027, 3404, 6487, -6339, -3619, 7977, 2, -7978, 3618, 6333, -6498, -3378, 8035, -284, -7906, 3890, 6129, -6691, -3070, 8094, -637, -7803, 4214, 5868, -6910, -2694, 8147, -1057, -7661, 4586, 5545, -7146, -2245, 8182, -1540, -7471, 4999, 5152, -7389, -1723, 8188, -2084, -7220, 5443, 4683, -7627, -1127, 8151, -2682, -6899, 5908, 4132, -7844, -456, 8056, -3327, -6495, 6378, 3493, -8023, 285, 7887, -4007, -5997, 6838, 2763, -8146, 1092, 7627, -4709, -5395, 7268, 1941, -8191, 1954, 7260, -5413, -4681, 7644, 1031, -8137, 2857, 6769, -6098, -3850, 7942, 40, -7962, 3783, 6142, -6738, -2901, 8133, -1020, -7642, 4706, 5368, -7301, -1839, 8189, -2128, -7159, 5597, 4442, -7755, -676, 8082, -3257, -6497, 6421, 3365, -8064, 569, 7784, -4375, -5645, 7137, 2148, -8190, 1868, 7272, -5440, -4600, 7700, 809, -8100, 3180, 6530, -6403, -3370, 8066, -619, -7761, 4460, 5550, -7212, -1974, 8190, -2095, -7150, 5649, 4337, -7810, -447, 8031, -3562, -6254, 6685, 2911, -8142, 1164, 7557, -4953, -5074, 7498, 1307, -8155, 2793, 6748, -6192, -3629, 8021, -419, -7810, 4363, 5603, -7198, -1961, 8190, -2191, -7079, 5782, 4142, -7888, -132, 7953, -3918, -5958, 6954, 2410, -8185, 1769, 7279, -5493, -4469, 7780, 482, -8028, 3635, 6160, -6800, -2666, 8170, -1540, -7377, 5341, 4622, -7726, -634, 8052, -3530, -6227, 6752, 2729, -8167, 1505, 7384, -5340, -4611, 7736, 585, -8041, 3602, 6162, -6817, -2606, 8176, -1668, -7305, 5488, 4431, -7810, -338, 7986, -3854, -5963, 6985, 2289, -8190, 2021, 7124, -5777, -4078, 7928, -110, -7871, 4270, 5610, -7241, -1776, 8180, -2563, -6821, 6184, 3534, -8064, 755, 7660, -4836, -5084, 7545, 1056, -8110, 3275, 6358, -6677, -2785, 8167, -1593, -7314, 5515, 4351, -7854, -131, 7923, -4134, -5698, 7202, 1813, -8181, 2602, 6774, -6264, -3388, 8096, -997, -7557, 5091, 4793, -7694, -616, 8027, -3749, -5989, 7008, 2170, -8191, 2295, 6937, -6084, -3614, 8058, -794, -7624, 4968, 4900, -7656, -702, 8039, -3715, -5999, 7012, 2139, -8191, 2371, 6882, -6168, -3479, 8087, -990, -7541, 5160, 4683, -7755, -388, 7968, -4034, -5730, 7215, 1719, -8171, 2826, 6596, -6502, -2973, 8158, -1580, -7277, 5644, 4120, -7950, 327, 7765, -4679, -5142, 7562, 897, -8066, 3635, 6021, -7023, -2069, 8187, -2545, -6752, 6354, 3164, -8142, 1436, 7328, -5583, -4168, 7943, -335, -7754, 4733, 5065, -7611, -740, 8030, -3831, -5850, 7162, 1766, -8170, 2895, 6515, -6619, -2733, 8180, -1950, -7065, 5996, 3626, -8077, 1008, 7496, -5316, -4441, 7869, -90, -7818, 4593, 5169, -7576, -798, 8034, -3846, -5812, 7206, 1640, -8157, 3085, 6366, -6779, -2433, 8190, -2327, -6838, 6303, 3168, -8149, 1579, 7227, -5796, -3846, 8040, -853, -7542, 5263, 4460, -7876, 153, 7784, -4720, -5015, 7663, 511, -7965, 4172, 5508, -7416, -1140, 8086, -3630, -5945, 7139, 1727, -8160, 3098, 6325, -6844, -2273, 8189, -2585, -6656, 6535, 2773, -8184, 2092, 6938, -6223, -3232, 8147, -1626, -7178, 5909, 3647, -8089, 1188, 7377, -5604, -4022, 8012, -782, -7544, 5308, 4355, -7926, 407, 7679, -5029, -4652, 7830, -68, -7789, 4766, 4910, -7733, -238, 7876, -4527, -5136, 7636, 508, -7945, 4310, 5328, -7546, -745, 7997, -4120, -5491, 7461, 944, -8038, 3955, 5623, -7389, -1111, 8066, -3822, -5729, 7326, 1241, -8088, 3715, 5807, -7280, -1339, 8101, -3641, -5863, 7247, 1400, -8110, 3596, 5891, -7231, -1429, 8112, -3584, -5897, 7230, 1422, -8111, 3601, 5878, -7246, -1383, 8103, -3651, -5836, 7277, 1308, -8092, 3729, 5767, -7325, -1200, 8072, -3840, -5674, 7385, 1056, -8046, 3979, 5553, -7458, -879, 8008, -4147, -5405, 7541, 665, -7959, 4341, 5225, -7633, -418, 7894, -4562, -5016, 7728, 134, -7813, 4805, 4771, -7826, 183, 7708, -5071, -4493, 7920, -536, -7580, 5352, 4176, -8009, 921, 7421, -5650, -3821, 8085, -1340, -7231, 5957, 3423, -8146, 1787, 7001, -6270, -2985, 8182, -2263, -6730, 6582, 2501) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L40C31_i
    );

    L40C32_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (134, 7798, 4877, -4667, -7874, -385, 7626, 5273, -4249, -7995, -868, 7440, 5624, -3847, -8082, -1313, 7244, 5932, -3463, -8140, -1721, 7044, 6202, -3102, -8174, -2091, 6847, 6435, -2767, -8190, -2423, 6655, 6635, -2459, -8190, -2718, 6473, 6804, -2181, -8181, -2977, 6305, 6947, -1933, -8164, -3201, 6152, 7065, -1718, -8144, -3390, 6018, 7161, -1535, -8123, -3547, 5905, 7236, -1386, -8103, -3670, 5814, 7293, -1271, -8086, -3762, 5746, 7334, -1189, -8073, -3823, 5701, 7358, -1142, -8066, -3853, 5682, 7366, -1129, -8065, -3852, 5688, 7360, -1151, -8070, -3820, 5718, 7338, -1206, -8081, -3758, 5773, 7301, -1296, -8096, -3665, 5852, 7246, -1420, -8115, -3540, 5953, 7173, -1578, -8136, -3382, 6076, 7081, -1768, -8157, -3191, 6218, 6966, -1992, -8176, -2965, 6378, 6828, -2247, -8188, -2705, 6553, 6662, -2532, -8191, -2408, 6740, 6467, -2847, -8181, -2074, 6935, 6239, -3189, -8154, -1702, 7134, 5976, -3556, -8105, -1293, 7332, 5673, -3945, -8029, -845, 7525, 5329, -4352, -7921, -361, 7706, 4940, -4772, -7774, 159, 7868, 4503, -5202, -7584, 713, 8006, 4018, -5633, -7345, 1299, 8110, 3481, -6060, -7051, 1911, 8174, 2894, -6475, -6697, 2545, 8189, 2255, -6869, -6278, 3194, 8146, 1568, -7232, -5791, 3851, 8037, 834, -7553, -5233, 4507, 7854, 58, -7821, -4601, 5150, 7588, -752, -8025, -3896, 5770, 7233, -1589, -8152, -3120, 6352, 6783, -2442, -8191, -2275, 6881, 6233, -3299, -8129, -1370, 7343, 5581, -4144, -7957, -413, 7720, 4828, -4962, -7663, 585, 7997, 3975, -5732, -7242, 1608, 8157, 3030, -6436, -6687, 2639, 8184, 2002, -7050, -5996, 3655, 8064, 904, -7554, -5172, 4634, 7786, -245, -7925, -4219, 5550, 7341, -1423, -8142, -3150, 6374, 6725, -2605, -8185, -1979, 7077, 5937, -3759, -8038, -729, 7631, 4984, -4854, -7689, 573, 8007, 3879, -5853, -7131, 1894, 8181, 2642, -6719, -6363, 3196, 8131, 1298, -7415, -5393, 4439, 7840, -118, -7906, -4236, 5575, 7301, -1564, -8161, -2917, 6561, 6513, -2993, -8153, -1470, 7349, 5486, -4353, -7864, 61, 7897, 4242, -5587, -7285, 1624, 8167, 2813, -6640, -6418, 3159, 8130, 1245, -7457, -5281, 4601, 7767, -407, -7988, -3903, 5883, 7072, -2075, -8190, -2330, 6937, 6057, -3687, -8036, -623, 7702, 4747, -5162, -7509, 1147, 8122, 3188, -6421, -6614, 2896, 8156, 1444, -7389, -5373, 4533, 7780, -405, -7996, -3833, 5965, 6991, -2268, -8191, -2061, 7102, 5808, -4040, -7939, -142, 7863, 4279, -5615, -7230, 1818, 8183, 2474, -6888, -6083, 3703, 8020, 489, -7765, -4544, 5393, 7357, -1560, -8170, -2694, 6769, 6212, -3542, -8052, -637, 7722, 4638, -5320, -7393, 1495, 8166, 2723, -6761, -6212, 3557, 8045, 585, -7745, -4569, 5396, 7341, -1628, -8177, -2565, 6863, 6078, -3753, -7999, -335, 7827, 4330, -5620, -7195, 1954, 8189, 2212, -7066, -5803, 4118, 7893, -116, -7953, -3913, 5972, 6933, -2468, -8181, -1663, 7342, 5364, -4640, -7701, 764, 8085, 3298, -6430, -6526, 3156, 8108, 905, -7656, -4736, 5288, 7377, -1606, -8179, -2474, 6946, 5932, -3995, -7920, 58, 7949, 3886, -6022, -6872, 2617, 8167, 1422, -7465, -5111, 4941, 7549, -1220, -8151, -2794, 6776, 6125, -3767, -7976, -148, 7903, 4021, -5935, -6927, 2546, 8171, 1444, -7467, -5087, 4986, 7516, -1328, -8163, -2641, 6880, 5981, -3979, -7911, 145, 7981, 3716, -6185, -6706, 2947, 8127, 972, -7660, -4661, 5416, 7266, -1925, -8191, -2007, 7229, 5470, -4610, -7678, 937, 8125, 2943, -6721, -6150, 3789, 7954, -4, -7957, -3779, 6162, 6704, -2983, -8119, -863, 7710, 4510, -5579, -7146, 2205, 8186, 1653, -7408, -5141, 4990, 7486, -1474, -8179, -2363, 7071, 5675, -4415, -7741, 796, 8112, 2990, -6719, -6122, 3867, 7922, -183, -8008, -3538, 6365, 6489, -3359, -8046, -366, 7876, 4005, -6027, -6788, 2896, 8122, 844, -7735, -4402, 5712, 7024, -2490, -8167, -1253, 7593, 4727, -5432, -7210, 2140, 8186, 1591, -7462, -4989, 5192, 7349, -1854, -8191, -1862, 7347, 5189, -4999, -7451, 1631, 8187, 2064, -7258, -5335, 4855, 7519, -1475, -8183, -2200, 7195, 5426, -4766, -7560, 1383, 8178, 2269, -7166, -5466, 4729, 7572, -1360, -8178, -2275, 7168, 5454, -4750, -7560, 1402, 8180, 2213, -7203, -5393, 4824, 7519, -1513, -8186, -2087, 7268, 5278, -4954, -7451, 1688, 8190, 1893, -7363, -5110, 5132, 7348, -1931, -8190, -1634, 7479, 4883, -5360, -7209, 2235, 8177, 1303, -7614, -4595, 5629, 7023, -2602, -8145, -906, 7755, 4238, -5936, -6787, 3025, 8083, 436, -7897, -3813, 6268, 6488, -3502, -7981, 102, 8024, 3310, -6619, -6121, 4022, 7825, -708, -8126, -2729, 6972, 5673, -4580, -7604, 1376, 8183, 2065, -7316, -5138, 5159, 7301, -2102, -8182, -1321, 7629, 4507, -5749, -6905, 2872, 8100, 496, -7895, -3776, 6327, 6399, -3677, -7922, 399, 8087, 2940, -6875, -5775, 4495, 7625, -1359, -8185, -2003, 7363, 5021, -5307, -7194, 2364, 8159, 967, -7766, -4134, 6081, 6609, -3394, -7989, 150, 8049, 3112, -6790, -5861, 4419, 7646, -1333, -8185, -1967, 7393, 4941, -5407, -7114, 2551, 8136, 708, -7854, -3851, 6314, 6372, -3772, -7877, 633, 8129, 2600, -7097, -5419, 4946, 7379, -2024, -8181, -1211, 7702, 4251, -6026, -6627, 3416, 7970, -284, -8083, -2889, 6950, 5611, -4754, -7471, 1834, 8187, 1359, -7658, -4343, 5968, 6662, -3381, -7975, 287, 8086, 2842, -6988, -5544, 4847, 7413, -1990, -8181, -1159, 7735, 4129, -6151, -6489, 3664, 7891, -647, -8139, -2462, 7199, 5205, -5218, -7192, 2484, 8134, 602, -7907, -3599, 6544, 6073, -4251, -7679, 1354, 8188, 1728, -7539, -4562, 5826, 6747, -3297, -7983, 309, 8098, 2715, -7086, -5358, 5090, 7251, -2394, -8142, -629, 7908, 3558, -6592, -5997, 4376, 7612, -1569, -8191, -1448, 7658, 4262, -6094, -6498, 3712, 7857, -838, -8164, -2144, 7381, 4834, -5622, -6881, 3120, 8014, -213, -8092, -2719, 7107, 5288, -5198, -7165, 2614, 8106, 302, -7998, -3176, 6858, 5634, -4841, -7367, 2206, 8155, 703, -7905, -3520, 6652, 5885, -4562, -7505, 1901, 8178, 992, -7828, -3758, 6501, 6049, -4372, -7588, 1703, 8186, 1168, -7778, -3893, 6415, 6135, -4273, -7627, 1614, 8188, 1233, -7761, -3929, 6397, 6145, -4271, -7623, 1636, 8187, 1187, -7779, -3866, 6449, 6081, -4363, -7578, 1766, 8182, 1030, -7831, -3703, 6568, 5939, -4549, -7486, 2006, 8166, 761, -7910, -3437, 6748, 5714, -4822, -7339, 2351, 8129, 378, -8003, -3062, 6977, 5396, -5175, -7124, 2798, 8056, -117, -8096, -2573, 7241, 4974, -5595, -6826, 3338, 7928, -724, -8167, -1966, 7520, 4436, -6065, -6425, 3960, 7720, -1437, -8191, -1235, 7788, 3770, -6563, -5903, 4646, 7409, -2248, -8137, -383, 8013, 2966, -7058, -5239, 5373, 6964, -3139, -7971, 586, 8158, 2020, -7514, -4417, 6107, 6360, -4086, -7658, 1656, 8182, 933, -7889, -3425, 6807, 5570, -5054, -7161, 2804, 8040, -284, -8130, -2260, 7423, 4577, -5997, -6446, 3990, 7686, -1605, -8184, -932, 7895, 3372, -6855, -5488, 5163, 7077, -2988, -7995, 534, 8158, 1963, -7559, -4273, 6254, 6179, -4374, -7511, 2091, 8145, 377, -8031, -2807, 7183, 4974, -5684, -6687, 3672, 7790, -1335, -8191, -1119, 7855, 3466, -6822, -5500, 5183, 7042, -3092, -7960, 731, 8176, 1687, -7679, -3954, 6513, 5871, -4787, -7278, 2651, 8054, -293, -8141, -2086, 7532, 4280, -6287, -6109, 4512, 7417, -2363, -8103, 20, 8108, 2318, -7441, -4460, 6159, 6227, -4374, -7481, 2233, 8118, 83, -8096, -2389, 7415, 4495, -6141, -6237, 4375, 7473, -2265, -8113, -21, 8106, 2299, -7462, -4392, 6231, 6134, -4518, -7396, 2456, 8079, -211, -8139, -2048, 7571, 4142, -6427, -5917, 4795, 7237, -2806, -8008, 608, 8174, 1629, -7730, -3740, 6709, 5567, -5196, -6979, 3302, 7874, -1171, -8191, -1041, 7910, 3171, -7058, -5068, 5697, 6594, -3933, -7647, 1891, 8150, 279, -8077, -2425, 7433, 4394, -6271, -6052, 4673, 7284, -2756, -8009, 652, 8180, 1490, -7791, -3527, 6870, 5316, -5487, -6744, 3735, 7711, -1740, -8162, -369, 8066, 2446, -7438, -4358, 6319, 5977, -4790, -7202, 2951, 7954, -927, -8191, -1153, 7898, 3152, -7101, -4947, 5853, 6420, -4239, -7486, 2360, 8077, -340, -8163, -1698, 7739, 3623, -6839, -5322, 5520, 6687, -3868, -7643, 1983, 8130, 15, -8128, -2009, 7635, 3875, -6690, -5507, 5348, 6807, -3696, -7704, 1830, 8146, 136, -8114, -2091, 7611, 3918, -6672, -5517, 5352, 6794, -3733, -7684, 1905, 8136, 23, -8131, -1947, 7671, 3755, -6788, -5351, 5531, 6647, -3976, -7578, 2206, 8091, -324, -8167, -1573, 7802, 3377, -7023, -4999, 5870, 6348, -4413, -7362, 2726, 7984, -903, -8191, -963, 7972, 2772, -7344, -4435, 6341, 5866, -5020, -6996, 3448, 7769, -1708, -8152, -113, 8126, 1922, -7700, -3632, 6894, 5157, -5755, -6428, 4338, 7382, -2718, -7979, 970, 8190, 817, -8013, -2562, 7456, 4178, -6552, -5596, 5342, 6747, -3891, -7585, 2263, 8069, -537, -8185, -1209, 7926, 2893, -7313, -4444, 6372, 5789, -5153, -6875, 3707, 7652, -2104, -8093, 413, 8179, 1289, -7912, -2932, 7303, 4442, -6387, -5760, 5201, 6828, -3801, -7607, 2244, 8065, -601, -8188, -1063, 7972, 2676, -7432, -4177, 6589, 5502, -5486, -6602, 4164, 7433, -2682, -7969, 1097, 8185, 524, -8083, -2120, 7664, 3627, -6953, -4992, 5975, 6159, -4774, -7089, 3395, 7747, -1896, -8115, 328, 8178, 1244, -7940, -2767, 7409, 4182, -6613, -5442, 5578, 6499, -4348, -7322, 2966, 7880, -1486, -8159, -44, 8151, 1564, -7860, -3027, 7297, 4378, -6488, -5577, 5460, 6581, -4252, -7361, 2905, 7891, -1467, -8159, -15, 8155, 1490, -7887, -2913, 7363, 4234, -6605, -5417, 5637, 6420, -4496, -7220, 3215, 7788, -1841, -8113, 414, 8185, 1020, -8008, -2418, 7586, 3736, -6938, -4938, 6084, 5987, -5054, -6857, 3878, 7519, -2594, -7963, 1238, 8172, 146, -8149, -1522, 7891, 2848, -7415, -4090, 6730, 5212, -5864, -6187, 4837, 6986, -3685, -7594, 2436, 7993, -1128, -8178, -207, 8144, 1528, -7897, -2806, 7444, 4004, -6801, -5096, 5985, 6051, -5022, -6850, 3934, 7472, -2754, -7908, 1509, 8144, -234, -8181, -1043, 8018, 2287, -7665, -3473, 7128, 4570, -6427, -5556, 5576, 6406, -4602, -7106, 3524, 7639, -2372, -7997, 1170, 8171, 52, -8165, -1268, 7975, 2450, -7614, -3574, 7087, 4614, -6412, -5552, 5601, 6367, -4678, -7045, 3659, 7572, -2571, -7942, 1433, 8146, -273, -8186, -888, 8059, 2025, -7775, -3118, 7337, 4143, -6761, -5084, 6054, 5921, -5237, -6644, 4324, 7236, -3335, -7692, 2288, 8001, -1205, -8165, 104, 8178, 991, -8047, -2065, 7771, 3096, -7363, -4069, 6826, 4964, -6177, -5772, 5423, 6477, -4585, -7070, 3672, 7542, -2705, -7889, 1697, 8104, -669, -8190, -366, 8143, 1388, -7970, -2385, 7672, 3337, -7260, -4235, 6737, 5062, -6118, -5811, 5408, 6468, -4625, -7028, 3777, 7481, -2882, -7826, 1948, 8057, -994, -8175, 30, 8178, 928, -8071, -1869, 7853, 2777, -7533, -3646, 7114, 4459, -6606, -5212, 6014, 5891, -5350, -6494, 4622, 7009, -3842, -7437, 3017, 7769, -2163, -8008, 1286, 8147, -401, -8191, -485, 8138, 1358, -7994, -2211, 7758, 3033, -7438, -3818, 7037, 4553, -6563, -5237, 6019, 5858, -5417, -6415, 4760, 6899, -4060, -7311, 3321, 7644, -2555, -7901, 1767, 8075, -969, -8172, 166, 8187, 632, -8127, -1421, 7989, 2188, -7780, -2933, 7500, 3643, -7156, -4318, 6750, 4948, -6290, -5533, 5777, 6065, -5221, -6544, 4624, 6963, -3995, -7324, 3337, 7621, -2658, -7858, 1962, 8030, -1259, -8141, 549, 8188, 158, -8176, -860, 8101, 1548, -7971, -2222, 7783, 2872, -7545, -3500, 7255, 4097, -6920, -4663, 6539, 5192, -6122, -5684, 5666, 6135, -5180, -6545, 4665, 6909, -4127, -7231, 3567, 7504, -2993, -7734, 2405, 7914, -1810, -8051, 1209, 8140, -608, -8186, 8, 8185, 585, -8144, -1171, 8059, 1744, -7937, -2305, 7774, 2847, -7577, -3372, 7344, 3874, -7081, -4356, 6786, 4810, -6466, -5241, 6118, 5643, -5750, -6018, 5359, 6363, -4952, -6679, 4528, 6964, -4092, -7220, 3643, 7444, -3187, -7640, 2722, 7803, -2254, -7939, 1782, 8043, -1311, -8121, 839, 8168, -371, -8190, -94, 8184, 551, -8154, -1003, 8098, 1444, -8021, -1878, 7919, 2299, -7799, -2710, 7656, 3107, -7497, -3492, 7318, 3861, -7125, -4218, 6915, 4557, -6693, -4883, 6457, 5191, -6211, -5485, 5953, 5761, -5688, -6023, 5413, 6267, -5133, -6496, 4845, 6707, -4555, -6905, 4258, 7085, -3961, -7251, 3660, 7401, -3359, -7537, 3056, 7658, -2755, -7767, 2453, 7860, -2155, -7942, 1857, 8010, -1564, -8068, 1272, 8112, -987, -8148, 703, 8171, -426, -8186, 152, 8190, 114, -8188, -377, 8175, 632, -8156, -882, 8129, 1125, -8096, -1363, 8056, 1592, -8012, -1817, 7961, 2032, -7907, -2243, 7848, 2446, -7786, -2643, 7719, 2831, -7652, -3015, 7580, 3189, -7508, -3359, 7433, 3521, -7358, -3677, 7281, 3825, -7205, -3969, 7126, 4104, -7050, -4235, 6973, 4358, -6898, -4477, 6822, 4588, -6749, -4695, 6676, 4794, -6606, -4890, 6537, 4979, -6471, -5064, 6406, 5142, -6345, -5217, 6285, 5285, -6230, -5351, 6175, 5409, -6126, -5465, 6078, 5515, -6035, -5562, 5994, 5602, -5958, -5640, 5923, 5673, -5894, -5702, 5867, 5726, -5846, -5748, 5827, 5764, -5813, -5778, 5801, 5785, -5795, -5791, 5792, 5791, -5794, -5789, 5797, 5781, -5807, -5772, 5819, 5756, -5836, -5738, 5856, 5714, -5881, -5689, 5908, 5657, -5940, -5622, 5975, 5582, -6014, -5539, 6056, 5490, -6102, -5438, 6150, 5380, -6203, -5319, 6257, 5252, -6315, -5181, 6375, 5103, -6439, -5023, 6503, 4935, -6572, -4844, 6640, 4745, -6713, -4642, 6785, 4532, -6860, -4419, 6935, 4297, -7012, -4171, 7088, 4037, -7166, -3898, 7242, 3751, -7320, -3600, 7395, 3440, -7471, -3276, 7544, 3102, -7617, -2924, 7685, 2737, -7754, -2546, 7817, 2345, -7878, -2139, 7934, 1925, -7988, -1706, 8034, 1478, -8077, -1245, 8113, 1004, -8144, -758, 8166, 504, -8183, -247, 8190, -19, -8190, 288, 8179, -564, -8161, 844, 8131, -1129, -8092, 1417, 8040, -1711, -7978, 2005, 7902, -2304, -7815, 2603, 7714, -2906, -7600, 3207, 7470, -3510, -7328, 3810, 7169, -4111, -6997, 4407, 6808, -4701, -6604, 4990, 6383, -5274, -6147, 5551, 5894, -5822, -5626, 6083, 5340, -6336, -5040, 6576, 4722, -6806, -4390, 7021, 4041, -7224, -3679, 7409, 3301, -7579, -2911, 7729, 2506, -7862, -2091, 7972, 1662, -8063, -1225, 8129, 777, -8173, -324, 8190, -139, -8183, 604, 8147, -1075, -8086, 1546, 7994, -2019, -7875, 2488, 7725, -2955, -7546, 3415, 7336, -3869, -7097, 4311, 6825, -4742, -6525, 5157, 6193, -5558, -5834, 5936, 5445, -6296, -5029, 6629, 4586, -6938, -4118, 7216, 3625, -7465, -3113, 7680, 2578, -7861, -2027, 8003, 1459, -8107, -880, 8170, 289, -8191, 307, 8168, -909, -8102, 1510, 7988, -2109, -7830, 2700, 7624, -3283, -7374, 3849, 7075, -4399, -6733, 4925, 6345, -5427, -5915, 5898, 5442, -6336, -4932, 6734, 4383, -7093, -3803, 7405, 3189, -7671, -2551, 7884, 1887, -8044, -1206, 8145, 510, -8190, 194, 8172, -904, -8094, 1611, 7952, -2312, -7748, 2999, 7480, -3669, -7151, 4313, 6760, -4928, -6312, 5504, 5805, -6040, -5248, 6526, 4638, -6961, -3986, 7335, 3292, -7649, -2565, 7893, 1807, -8067, -1029, 8166, 234, -8190, 567, 8133, -1370, -7998, 2163, 7782, -2941, -7488, 3694, 7114, -4415, -6666, 5094, 6144, -5726, -5555, 6298, 4902, -6809, -4192, 7247, 3430, -7609, -2627, 7886, 1787, -8078, -924, 8176, 42, -8182, 844, 8089, -1727, -7901, 2593, 7614, -3435, -7235, 4237, 6762, -4994, -6203, 5690, 5560, -6320, -4844, 6870, 4059, -7336, -3218, 7705, 2327, -7976, -1402, 8138, 450, -8191, 511, 8130, -1473, -7956, 2418, 7667, -3335, -7268, 4208, 6760, -5026, -6152, 5773, 5447, -6439, -4659, 7011, 3793, -7481, -2868, 7836, 1890, -8073, -880, 8182, -152, -8164, 1184, 8013, -2205, -7732, 3194, 7321, -4137, -6789, 5013, 6137, -5812, -5381, 6514, 4526, -7110, -3591, 7583, 2586, -7927, -1533, 8130, 445, -8191, 655, 8101, -1750, -7865, 2817, 7481, -3838, -6957, 4791, 6298, -5659, -5517, 6422, 4625, -7066, -3640, 7574, 2578, -7937, -1462, 8142, 309, -8187, 854, 8064, -2007, -7778, 3122, 7328, -4179, -6725, 5152, 5975, -6023, -5098, 6767, 4105, -7371, -3021, 7815, 1864, -8093, -663, 8190, -560, -8107, 1775, 7840, -2956, -7395, 4074, 6776, -5104, -6000, 6018, 5078, -6798, -4035, 7418, 2889, -7866, -1671, 8124, 406, -8188, 873, 8050, -2138, -7715, 3353, 7184, -4492, -6472, 5520, 5591, -6414, -4566, 7145, 3417, -7696, -2176, 8047, 871, -8189, 461, 8113, -1788, -7821, 3070, 7315, -4276, -6610, 5368, 5719, -6319, -4668, 7096, 3481, -7680, -2194, 8048, 837, -8190, 547, 8096, -1923, -7770, 3247, 7214, -4482, -6447, 5589, 5483, -6536, -4355, 7289, 3089, -7827, -1727, 8127, 304, -8181, 1131, 7981, -2538, -7534, 3869, 6847, -5086, -5943, 6144, 4845, -7012, -3589, 7655, 2210, -8055, -757, 8190, -729, -8059, 2194, 7658, -3593, -7002, 4876, 6105, -6000, -5000, 6922, 3719, -7612, -2307, 8040, 808, -8191, 723, 8055, -2236, -7635, 3672, 6941, -4985, -5998, 6122, 4834, -7043, -3492, 7709, 2015, -8096, -461, 8184, -1117, -7969, 2657, 7453, -4104, -6656, 5399, 5602, -6495, -4332, 7343, 2888, -7912, -1330, 8174, -288, -8118, 1898, 7739, -3440, -7054, 4848, 6083, -6068, -4865, 7046, 3445, -7742, -1881, 8121, 232, -8169, 1429, 7877, -3038, -7257, 4523, 6327, -5825, -5129, 6881, 3707, -7649, -2123, 8088, 441, -8181, 1264, 7916, -2921, -7305, 4453, 6367, -5795, -5146, 6881, 3689, -7663, -2064, 8101, 338, -8174, 1407, 7872, -3094, -7209, 4643, 6208, -5982, -4917, 7044, 3390, -7781, -1701, 8150, -77, -8134, 1854, 7727, -3550, -6948, 5077, 5828, -6364, -4423, 7341, 2794, -7963, -1025, 8190, -802, -8012, 2593, 7429, -4261, -6473, 5716, 5184, -6887, -3628, 7707, 1880, -8135, -31, 8141, -1826, -7724, 3592, 6900, -5176, -5712, 6489, 4216, -7463, -2493, 8038, 629, -8185, 1272, 7888, -3112, -7162, 4785, 6041, -6202, -4586, 7279, 2871, -7957, -993, 8190, -947, -7967, 2838, 7291, -4575, -6201, 6054, 4752, -7193, -3028, 7919, 1122, -8190, 852, 7983, -2783, -7310, 4555, 6203, -6064, -4727, 7216, 2964, -7941, -1021, 8190, -991, -7948, 2946, 7220, -4730, -6052, 6227, 4507, -7346, -2683, 8013, 685, -8184, 1359, 7843, -3325, -7010, 5085, 5729, -6529, -4083, 7559, 2170, -8110, -115, 8138, -1955, -7641, 3902, 6644, -5601, -5212, 6935, 3431, -7817, -1421, 8182, -691, -8005, 2760, 7289, -4650, -6083, 6230, 4460, -7394, -2531, 8054, 423, -8166, 1717, 7713, -3747, -6728, 5519, 5269, -6913, -3441, 7823, 1364, -8187, 812, 7969, -2938, -7186, 4858, 5884, -6436, -4158, 7552, 2125, -8125, 65, 8106, -2257, -7496, 4288, 6332, -6009, -4698, 7287, 2710, -8028, -517, 8168, -1723, -7696, 3836, 6640, -5665, -5079, 7066, 3125, -7932, -929, 8188, -1346, -7814, 3521, 6832, -5428, -5316, 6914, 3379, -7862, -1173, 8190, -1133, -7872, 3353, 6924, -5311, -5422, 6847, 3478, -7835, -1250, 8190, -1086, -7881, 3337, 6925, -5321, -5400, 6870, 3424, -7857, -1162, 8190, -1204, -7843, 3473, 6835, -5457, -5251, 6983, 3217, -7922, -907, 8185, -1488, -7751, 3758, 6646, -5712, -4967, 7173, 2851, -8016, -484, 8158, -1933, -7586, 4183, 6342, -6070, -4535, 7421, 2319, -8115, 108, 8081, -2532, -7322, 4731, 5898, -6508, -3937, 7695, 1611, -8183, 866, 7919, -3270, -6926, 5376, 5288, -6989, -3156, 7952, 723, -8174, 1781, 7626, -4124, -6359, 6081, 4484, -7465, -2179, 8137, -340, -8033, 2831, 7153, -5055, -5580, 6792, 3461, -7874, -1002, 8186, -1563, -7696, 3977, 6445, -6006, -4556, 7440, 2207, -8138, 365, 8021, -2908, -7100, 5161, 5458, -6899, -3261, 7937, 727, -8170, 1886, 7565, -4312, -6183, 6296, 4157, -7635, -1698, 8182, -945, -7877, 3492, 6745, -5680, -4903, 7271, 2537, -8098, 101, 8063, -2735, -7170, 5080, 5505, -6886, -3246, 7951, 630, -8159, 2058, 7479, -4529, -5983, 6507, 3827, -7777, -1247, 8190, -1478, -7699, 4042, 6349, -6163, -4290, 7597, 1745, -8183, 1000, 7846, -3638, -6622, 5868, 4642, -7436, -2130, 8155, -632, -7942, 3324, 6812, -5641, -4894, 7306, 2402, -8126, 373, 7998, -3111, -6933, 5487, 5049, -7222, -2566, 8104, -227, -8026, 2997, 6989, -5416, -5115, 7187, 2621, -8098, 192, 8030, -2989, -6989, 5426, 5092, -7207, -2572, 8107, -271, -8012, 3084, 6927, -5523, -4983, 7278, 2413, -8131, 461, 7967, -3284, -6803, 5697, 4779, -7397, -2147, 8160, -763, -7889, 3580, 6607, -5946, -4479, 7550, 1768, -8186, 1174, 7762, -3971, -6331, 6255, 4071, -7727, -1275, 8188, -1694, -7574, 4444, 5957, -6612, -3550, 7905, 665, -8149, 2313, 7301, -4987, -5474, 6994, 2904, -8063, 60, 8039, -3024, -6924, 5579, 4861, -7378, -2131, 8166, -898, -7834, 3808, 6417, -6197, -4109, 7727, 1224, -8186, 1835, 7498, -4644, -5758, 6803, 3202, -8007, -192, 8078, -2854, -7002, 5496, 4925, -7359, -2140, 8168, -958, -7806, 3921, 6314, -6325, -3906, 7812, 925, -8166, 2195, 7325, -5000, -5410, 7073, 2694, -8109, 422, 7945, -3483, -6603, 6030, 4274, -7682, -1303, 8185, -1869, -7461, 4764, 5609, -6946, -2908, 8077, -242, -7983, 3358, 6670, -5967, -4335, 7664, 1329, -8187, 1886, 7444, -4815, -5549, 7001, 2786, -8102, 414, 7937, -3556, -6529, 6142, 4091, -7768, -1005, 8166, -2247, -7272, 5145, 5217, -7230, -2328, 8160, -940, -7784, 4061, 6152, -6533, -3527, 7951, 323, -8082, 2936, 6896, -5723, -4583, 7576, 1513, -8190, 1809, 7454, -4839, -5487, 7071, 2606, -8134, 712, 7842, -3918, -6240, 6471, 3588, -7943, -330, 8077, -2991, -6848, 5809, 4453, -7646, -1299, 8181, -2083, -7320, 5112, 5201, -7269, -2185, 8175, -1214, -7671, 4406, 5834, -6840, -2981, 8083, -399, -7917, 3712, 6361, -6380, -3685, 7926, 353, -8075, 3045, 6791, -5909, -4299, 7723, 1034, -8161, 2419, 7135, -5444, -4826, 7492, 1642, -8191, 1843, 7405, -5000, -5273, 7249, 2175, -8180, 1324, 7611, -4587, -5645, 7008, 2634, -8141, 867, 7766, -4215, -5950, 6781, 3021, -8087, 476, 7880, -3890, -6194, 6576, 3338, -8027, 151, 7960, -3618, -6384, 6401, 3589, -7970, -106, 8014, -3404, -6524, 6263, 3775, -7921, -295, 8050, -3248, -6620, 6165, 3899, -7887, -417, 8069, -3154, -6674, 6110, 3963, -7869, -470, 8077, -3123, -6688, 6100, 3968, -7871, -456, 8073, -3154, -6663, 6135, 3913, -7891, -373, 8057, -3248, -6597, 6215, 3797, -7927, -223, 8026, -3403, -6489, 6336, 3620, -7977, -5, 7978, -3617, -6336, 6496, 3379, -8035, 281, 7906, -3889, -6131, 6689, 3072, -8095, 634, 7803, -4213, -5871, 6908, 2695, -8148, 1053, 7661, -4585, -5548, 7144, 2247, -8183, 1537, 7470, -4998, -5155, 7387, 1725, -8189, 2081, 7220, -5442, -4686, 7625, 1128, -8153, 2679, 6899, -5907, -4135, 7842, 457, -8058, 3324, 6495, -6378, -3496, 8022, -284, -7889, 4004, 5997, -6838, -2766, 8145, -1091, -7629, 4706, 5396, -7268, -1944, 8190, -1953, -7262, 5410, 4682, -7644, -1034, 8137, -2856, -6772, 6095, 3851, -7942, -43, 7961, -3782, -6145, 6735, 2902, -8134, 1016, 7642, -4705, -5371, 7299, 1840, -8190, 2124, 7159, -5597, -4445, 7753, 677, -8083, 3254, 6497, -6420, -3369, 8062, -568, -7786, 4372, 5645, -7136, -2151, 8189, -1866, -7274, 5437, 4601, -7700, -813, 8099, -3179, -6533, 6401, 3371, -8067, 616, 7761, -4459, -5553, 7210, 1976, -8191, 2091, 7150, -5648, -4341, 7808, 448, -8033, 3558, 6255, -6684, -2914, 8140, -1162, -7559, 4950, 5075, -7498, -1310, 8155, -2792, -6751, 6190, 3630, -8021, 415, 7810, -4362, -5606, 7196, 1962, -8191, 2188, 7080, -5781, -4145, 7886, 134, -7955, 3915, 5959, -6953, -2414, 8184, -1767, -7281, 5490, 4471, -7780, -486, 8027, -3634, -6163, 6798, 2667, -8171, 1537, 7377, -5340, -4625, 7725, 636, -8054, 3527, 6228, -6751, -2732, 8166, -1504, -7386, 5337, 4612, -7736, -588, 8041, -3601, -6165, 6815, 2607, -8177, 1664, 7305, -5487, -4434, 7808, 340, -7987, 3850, 5964, -6985, -2292, 8189, -2020, -7126, 5774, 4079, -7928, 106, 7870, -4268, -5613, 7238, 1778, -8181, 2560, 6821, -6183, -3537, 8062, -753, -7662, 4833, 5085, -7545, -1060, 8110, -3274, -6361, 6674, 2787, -8168, 1589, 7314, -5514, -4355, 7852, 133, -7924, 4131, 5698, -7202, -1817, 8180, -2600, -6777, 6261, 3389, -8096, 993, 7557, -5090, -4797, 7692, 618, -8029, 3746, 5989, -7007, -2174, 8190, -2294, -6940, 6081, 3616, -8059, 791, 7624, -4967, -4904, 7654, 703, -8041, 3712, 6000, -7012, -2143, 8190, -2370, -6884, 6165, 3481, -8088, 987, 7541, -5159, -4687, 7753, 389, -7969, 4030, 5731, -7214, -1722, 8170, -2825, -6599, 6499, 2975, -8159, 1577, 7277, -5643, -4124, 7948, -326, -7766, 4676, 5144, -7562, -901, 8066, -3633, -6024, 7020, 2071, -8188, 2542, 6753, -6353, -3168, 8140, -1434, -7330, 5580, 4170, -7943, 331, 7754, -4732, -5068, 7609, 742, -8032, 3828, 5851, -7162, -1770, 8170, -2894, -6518, 6616, 2734, -8181, 1946, 7065, -5995, -3629, 8075, -1007, -7498, 5313, 4442, -7869, 86, 7818, -4592, -5172, 7573, 799, -8036, 3842, 5813, -7206, -1644, 8156, -3083, -6369, 6776, 2435, -8191, 2323, 6839, -6303, -3172, 8148, -1577, -7229, 5793, 3847, -8040, 849, 7542, -5262, -4463, 7874, -151, -7786, 4717, 5016, -7663, -515, 7964, -4170, -5511, 7414, 1142, -8088, 3626, 5946, -7138, -1731, 8159, -3096, -6328, 6841, 2274, -8190, 2581, 6657, -6534, -2777, 8183, -2090, -6940, 6220, 3234, -8148, 1623, 7178, -5908, -3651, 8088, -1186, -7379, 5601, 4024, -8013, 778, 7544, -5307, -4359, 7924, -405, -7681, 5026, 4654, -7830, 64, 7789, -4765, -4914, 7731, 240, -7877, 4524, 5138, -7636, -512, 7945, -4308, -5331, 7544, 747, -7998, 4116, 5492, -7461, -948, 8037, -3954, -5626, 7386, 1113, -8068, 3818, 5730, -7326, -1245, 8087, -3714, -5811, 7278, 1341, -8102, 3637, 5864, -7246, -1404, 8109, -3594, -5894, 7229, 1431, -8113, 3580, 5899, -7229, -1426, 8111, -3599, -5881, 7244, 1385, -8105, 3647, 5837, -7277, -1312, 8091, -3728, -5770, 7322, 1202, -8073, 3836, 5676, -7384, -1060, 8045, -3977, -5556, 7456, 881, -8009, 4144, 5406, -7540, -669, 7959, -4339, -5229, 7631, 420, -7896, 4559, 5018, -7728, -138, 7813, -4803, -4775, 7824, -181, -7710, 5067, 4495, -7920, 532, 7581, -5351, -4179, 8008, -919, -7424, 5647, 3822, -8086, 1336, 7231, -5955, -3427, 8144, -1785, -7003, 6267, 2987, -8182, 2259, 6731, -6581, -2505) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L40C32_i
    );

    L40C33_instance: entity work.LHM_ALL
    generic map(
     rom_cos => (-131, -7798, -4880, 4663, 7873, 387, -7626, -5276, 4246, 7995, 870, -7439, -5627, 3843, 8081, 1315, -7243, -5936, 3459, 8139, 1723, -7044, -6205, 3098, 8173, 2093, -6846, -6438, 2763, 8189, 2425, -6654, -6637, 2455, 8189, 2720, -6472, -6807, 2176, 8180, 2979, -6304, -6950, 1929, 8163, 3203, -6151, -7067, 1714, 8143, 3392, -6017, -7163, 1531, 8121, 3548, -5904, -7239, 1382, 8101, 3672, -5812, -7296, 1267, 8084, 3764, -5744, -7336, 1185, 8072, 3824, -5700, -7360, 1138, 8065, 3854, -5681, -7369, 1125, 8064, 3854, -5687, -7362, 1147, 8069, 3822, -5717, -7341, 1202, 8079, 3760, -5772, -7303, 1292, 8095, 3667, -5851, -7249, 1416, 8114, 3542, -5952, -7176, 1574, 8135, 3384, -6075, -7083, 1764, 8156, 3193, -6217, -6969, 1988, 8174, 2967, -6377, -6830, 2243, 8187, 2707, -6552, -6665, 2529, 8190, 2410, -6739, -6470, 2843, 8181, 2076, -6934, -6242, 3186, 8154, 1704, -7133, -5979, 3553, 8105, 1295, -7332, -5677, 3941, 8029, 847, -7525, -5332, 4348, 7920, 363, -7706, -4943, 4769, 7774, -157, -7868, -4507, 5198, 7584, -711, -8006, -4021, 5630, 7345, -1297, -8111, -3485, 6057, 7051, -1909, -8175, -2898, 6472, 6698, -2543, -8190, -2259, 6866, 6279, -3192, -8148, -1571, 7229, 5792, -3850, -8039, -838, 7551, 5234, -4505, -7856, -62, 7819, 4602, -5149, -7590, 748, 8023, 3898, -5769, -7235, 1585, 8151, 3121, -6351, -6785, 2438, 8190, 2277, -6881, -6236, 3295, 8129, 1372, -7343, -5584, 4141, 7956, 414, -7720, -4831, 4958, 7664, -583, -7998, -3979, 5729, 7242, -1607, -8158, -3034, 6433, 6687, -2637, -8185, -2005, 7048, 5997, -3654, -8066, -908, 7552, 5173, -4633, -7788, 241, 7923, 4221, -5549, -7343, 1420, 8141, 3151, -6373, -6727, 2601, 8184, 1981, -7077, -5940, 3756, 8038, 731, -7631, -4988, 4851, 7689, -571, -8008, -3883, 5850, 7131, -1892, -8182, -2645, 6716, 6364, -3195, -8132, -1301, 7413, 5394, -4437, -7842, 114, 7905, 4237, -5574, -7303, 1560, 8160, 2918, -6560, -6516, 2990, 8152, 1471, -7349, -5489, 4349, 7864, -59, -7897, -4245, 5584, 7285, -1622, -8168, -2817, 6638, 6419, -3157, -8131, -1249, 7455, 5282, -4600, -7769, 403, 7986, 3904, -5882, -7075, 2072, 8189, 2332, -6937, -6059, 3683, 8035, 624, -7702, -4750, 5159, 7509, -1146, -8122, -3192, 6419, 6614, -2895, -8157, -1448, 7386, 5374, -4532, -7782, 402, 7995, 3835, -5964, -6993, 2264, 8190, 2062, -7102, -5811, 4037, 7938, 144, -7864, -4282, 5612, 7230, -1816, -8184, -2477, 6886, 6083, -3702, -8021, -492, 7763, 4546, -5392, -7359, 1556, 8169, 2695, -6768, -6215, 3538, 8052, 639, -7722, -4642, 5317, 7393, -1494, -8167, -2726, 6759, 6213, -3556, -8046, -589, 7743, 4570, -5395, -7343, 1625, 8176, 2566, -6862, -6081, 3750, 7998, 337, -7827, -4333, 5617, 7195, -1952, -8190, -2216, 7063, 5804, -4117, -7895, 113, 7951, 3914, -5971, -6935, 2465, 8180, 1664, -7342, -5367, 4637, 7701, -763, -8086, -3302, 6427, 6527, -3154, -8109, -908, 7654, 4737, -5287, -7379, 1602, 8178, 2475, -6946, -5935, 3992, 7920, -57, -7949, -3889, 6019, 6872, -2616, -8168, -1425, 7463, 5112, -4940, -7551, 1217, 8150, 2795, -6775, -6128, 3764, 7976, 150, -7903, -4024, 5932, 6927, -2545, -8172, -1448, 7465, 5088, -4985, -7518, 1325, 8162, 2643, -6879, -5984, 3976, 7911, -144, -7981, -3719, 6183, 6706, -2945, -8128, -975, 7658, 4662, -5415, -7268, 1922, 8190, 2008, -7228, -5473, 4607, 7678, -935, -8126, -2946, 6719, 6151, -3788, -7956, 1, 7956, 3780, -6161, -6706, 2980, 8118, 865, -7710, -4512, 5576, 7146, -2204, -8187, -1656, 7406, 5142, -4989, -7488, 1471, 8178, 2364, -7070, -5677, 4412, 7741, -795, -8113, -2993, 6717, 6123, -3865, -7923, 179, 8006, 3539, -6365, -6492, 3355, 8045, 367, -7877, -4009, 6025, 6788, -2895, -8124, -847, 7734, 4403, -5711, -7026, 2487, 8166, 1255, -7593, -4730, 5430, 7210, -2139, -8187, -1594, 7460, 4990, -5191, -7351, 1851, 8190, 1863, -7347, -5192, 4996, 7451, -1629, -8188, -2067, 7256, 5336, -4854, -7521, 1471, 8182, 2201, -7195, -5428, 4763, 7560, -1382, -8179, -2272, 7164, 5467, -4728, -7574, 1357, 8177, 2276, -7167, -5457, 4747, 7560, -1401, -8181, -2216, 7201, 5394, -4823, -7521, 1510, 8185, 2089, -7268, -5281, 4951, 7451, -1687, -8191, -1897, 7361, 5111, -5132, -7350, 1928, 8189, 1635, -7479, -4885, 5358, 7209, -2234, -8178, -1307, 7612, 4596, -5629, -7025, 2599, 8145, 907, -7756, -4241, 5933, 6787, -3024, -8084, -439, 7896, 3814, -6268, -6490, 3499, 7981, -101, -8025, -3313, 6617, 6121, -4021, -7827, 705, 8125, 2730, -6972, -5675, 4577, 7604, -1375, -8184, -2068, 7314, 5139, -5159, -7303, 2099, 8181, 1322, -7629, -4509, 5747, 6905, -2871, -8101, -500, 7893, 3777, -6327, -6401, 3674, 7922, -398, -8088, -2943, 6873, 5776, -4494, -7627, 1356, 8184, 2004, -7363, -5023, 5304, 7194, -2363, -8161, -970, 7764, 4135, -6081, -6611, 3392, 7989, -149, -8050, -3115, 6788, 5862, -4418, -7648, 1330, 8184, 1968, -7393, -4943, 5405, 7114, -2550, -8138, -711, 7852, 3852, -6313, -6375, 3769, 7877, -632, -8129, -2603, 7095, 5419, -4946, -7381, 2021, 8180, 1212, -7702, -4254, 6024, 6627, -3415, -7972, 281, 8082, 2890, -6950, -5613, 4752, 7471, -1833, -8188, -1362, 7657, 4343, -5968, -6664, 3378, 7975, -286, -8087, -2845, 6986, 5544, -4846, -7415, 1987, 8180, 1160, -7735, -4132, 6149, 6489, -3663, -7892, 644, 8138, 2462, -7200, -5208, 5216, 7191, -2483, -8136, -605, 7906, 3599, -6544, -6075, 4248, 7678, -1353, -8189, -1731, 7538, 4563, -5825, -6749, 3295, 7983, -309, -8099, -2717, 7084, 5358, -5090, -7253, 2392, 8141, 629, -7909, -3561, 6590, 5997, -4375, -7614, 1566, 8190, 1449, -7658, -4264, 6092, 6499, -3711, -7859, 835, 8163, 2145, -7382, -4837, 5619, 6881, -3119, -8015, 210, 8090, 2720, -7107, -5290, 5196, 7165, -2614, -8107, -305, 7997, 3176, -6858, -5636, 4838, 7367, -2205, -8156, -706, 7904, 3521, -6652, -5887, 4560, 7504, -1900, -8179, -995, 7826, 3758, -6501, -6051, 4369, 7588, -1702, -8187, -1171, 7776, 3894, -6415, -6137, 4271, 7626, -1614, -8189, -1236, 7759, 3929, -6397, -6147, 4268, 7623, -1635, -8188, -1190, 7778, 3867, -6449, -6083, 4361, 7578, -1766, -8183, -1033, 7830, 3704, -6568, -5941, 4546, 7486, -2005, -8167, -763, 7908, 3437, -6748, -5716, 4820, 7339, -2351, -8130, -381, 8002, 3063, -6977, -5398, 5173, 7124, -2797, -8057, 114, 8095, 2574, -7242, -4976, 5593, 6826, -3338, -7929, 721, 8166, 1966, -7520, -4438, 6063, 6425, -3960, -7722, 1435, 8190, 1236, -7788, -3772, 6561, 5903, -4646, -7410, 2245, 8136, 384, -8013, -2969, 7056, 5239, -5372, -6966, 3137, 7971, -585, -8159, -2023, 7513, 4417, -6107, -6362, 4084, 7658, -1656, -8183, -935, 7887, 3426, -6807, -5572, 5052, 7160, -2803, -8041, 282, 8129, 2261, -7423, -4579, 5995, 6446, -3990, -7687, 1602, 8184, 932, -7896, -3375, 6853, 5488, -5163, -7078, 2986, 7995, -533, -8159, -1966, 7558, 4274, -6254, -6181, 4372, 7510, -2091, -8146, -379, 8030, 2808, -7183, -4976, 5682, 6687, -3671, -7791, 1332, 8190, 1120, -7856, -3468, 6820, 5501, -5183, -7043, 3090, 7960, -731, -8177, -1689, 7677, 3954, -6513, -5873, 4785, 7278, -2650, -8056, 291, 8140, 2086, -7532, -4282, 6285, 6109, -4512, -7419, 2361, 8102, -20, -8109, -2320, 7440, 4460, -6159, -6229, 4372, 7480, -2233, -8119, -86, 8094, 2390, -7416, -4497, 6139, 6236, -4375, -7474, 2263, 8112, 22, -8107, -2301, 7460, 4392, -6231, -6136, 4516, 7396, -2456, -8080, 208, 8138, 2048, -7571, -4144, 6425, 5917, -4795, -7238, 2803, 8008, -607, -8175, -1631, 7729, 3740, -6710, -5569, 5194, 6979, -3301, -7875, 1169, 8190, 1041, -7910, -3173, 7056, 5068, -5697, -6596, 3931, 7646, -1891, -8151, -281, 8076, 2425, -7433, -4396, 6269, 6052, -4673, -7285, 2754, 8009, -651, -8180, -1493, 7789, 3527, -6870, -5318, 5485, 6743, -3735, -7713, 1737, 8161, 370, -8067, -2449, 7437, 4358, -6319, -5979, 4788, 7202, -2951, -7955, 925, 8190, 1153, -7898, -3154, 7100, 4947, -5853, -6422, 4237, 7486, -2360, -8078, 338, 8162, 1698, -7740, -3625, 6838, 5322, -5520, -6689, 3865, 7642, -1982, -8132, -18, 8127, 2009, -7636, -3877, 6688, 5507, -5348, -6809, 3694, 7704, -1830, -8147, -139, 8113, 2092, -7611, -3920, 6670, 5517, -5352, -6796, 3731, 7683, -1905, -8137, -26, 8130, 1947, -7671, -3757, 6786, 5351, -5531, -6649, 3974, 7577, -2206, -8092, 322, 8166, 1573, -7803, -3379, 7021, 4999, -5871, -6350, 4411, 7361, -2726, -7986, 901, 8190, 963, -7973, -2774, 7343, 4435, -6342, -5867, 5018, 6996, -3448, -7770, 1706, 8151, 114, -8127, -1924, 7699, 3632, -6894, -5159, 5754, 6428, -4338, -7383, 2716, 7978, -970, -8191, -819, 8012, 2562, -7456, -4180, 6550, 5596, -5343, -6749, 3889, 7584, -2262, -8070, 535, 8183, 1209, -7927, -2895, 7312, 4444, -6373, -5791, 5151, 6874, -3707, -7653, 2102, 8092, -413, -8180, -1291, 7910, 2932, -7304, -4444, 6385, 5760, -5201, -6829, 3799, 7607, -2244, -8066, 599, 8187, 1063, -7973, -2678, 7430, 4177, -6590, -5503, 5484, 6602, -4164, -7435, 2680, 7968, -1097, -8186, -526, 8082, 2120, -7665, -3629, 6951, 4992, -5975, -6160, 4773, 7089, -3396, -7749, 1894, 8114, -328, -8178, -1246, 7938, 2767, -7410, -4184, 6611, 5441, -5578, -6501, 4347, 7321, -2966, -7881, 1484, 8159, 44, -8151, -1566, 7859, 3027, -7298, -4380, 6487, 5577, -5460, -6583, 4251, 7361, -2905, -7892, 1465, 8158, 15, -8156, -1492, 7886, 2912, -7363, -4236, 6603, 5416, -5637, -6422, 4494, 7219, -3215, -7789, 1839, 8112, -414, -8186, -1021, 8006, 2418, -7586, -3738, 6937, 4938, -6084, -5989, 5053, 6856, -3878, -7521, 2592, 7962, -1239, -8173, -147, 8147, 1522, -7892, -2850, 7413, 4090, -6731, -5214, 5862, 6186, -4838, -6988, 3683, 7594, -2436, -7994, 1126, 8178, 207, -8145, -1530, 7896, 2806, -7444, -4006, 6800, 5096, -5985, -6052, 5020, 6850, -3934, -7474, 2752, 7907, -1509, -8145, 232, 8180, 1043, -8019, -2289, 7664, 3473, -7129, -4572, 6426, 5556, -5577, -6408, 4600, 7106, -3524, -7640, 2370, 7996, -1170, -8172, -53, 8164, 1268, -7976, -2451, 7613, 3574, -7088, -4616, 6411, 5552, -5602, -6368, 4676, 7045, -3659, -7573, 2569, 7941, -1433, -8147, 272, 8185, 888, -8060, -2027, 7774, 3118, -7338, -4144, 6759, 5084, -6055, -5923, 5236, 6643, -4324, -7237, 3333, 7691, -2288, -8003, 1203, 8164, -104, -8179, -993, 8046, 2065, -7772, -3097, 7361, 4068, -6827, -4966, 6175, 5772, -5424, -6478, 4583, 7070, -3672, -7543, 2703, 7888, -1698, -8105, 668, 8189, 366, -8144, -1390, 7969, 2384, -7673, -3339, 7259, 4235, -6738, -5064, 6116, 5810, -5409, -6469, 4624, 7027, -3778, -7482, 2880, 7826, -1948, -8058, 992, 8175, -30, -8179, -929, 8070, 1868, -7854, -2779, 7532, 3645, -7114, -4460, 6605, 5211, -6014, -5892, 5349, 6493, -4622, -7010, 3840, 7436, -3018, -7770, 2161, 8007, -1286, -8148, 400, 8190, 484, -8139, -1359, 7993, 2211, -7759, -3034, 7437, 3817, -7037, -4555, 6561, 5236, -6020, -5859, 5415, 6414, -4760, -6900, 4058, 7310, -3321, -7646, 2554, 7900, -1768, -8076, 968, 8171, -166, -8188, -634, 8126, 1420, -7990, -2190, 7779, 2932, -7501, -3645, 7155, 4318, -6751, -4950, 6289, 5533, -5778, -6066, 5220, 6543, -4625, -6964, 3994, 7323, -3337, -7623, 2657, 7858, -1963, -8032, 1257, 8141, -549, -8189, -160, 8175, 859, -8102, -1550, 7970, 2221, -7784, -2874, 7544, 3499, -7255, -4098, 6918, 4662, -6540, -5193, 6120, 5684, -5667, -6136, 5179, 6544, -4665, -6910, 4126, 7230, -3568, -7505, 2992, 7733, -2406, -7916, 1809, 8050, -1210, -8141, 607, 8185, -9, -8186, -586, 8143, 1171, -8060, -1746, 7936, 2304, -7775, -2848, 7576, 3371, -7345, -3876, 7080, 4355, -6787, -4812, 6465, 5240, -6119, -5644, 5749, 6017, -5360, -6364, 4951, 6678, -4529, -6965, 4091, 7220, -3643, -7445, 3185, 7639, -2722, -7804, 2253, 7938, -1783, -8044, 1310, 8120, -839, -8169, 370, 8189, 93, -8185, -552, 8153, 1002, -8099, -1446, 8020, 1877, -7920, -2300, 7798, 2710, -7657, -3108, 7496, 3491, -7319, -3863, 7124, 4217, -6916, -4558, 6692, 4882, -6458, -5193, 6210, 5485, -5954, -5763, 5687, 6022, -5414, -6268, 5132, 6495, -4846, -6709, 4554, 6904, -4259, -7086, 3960, 7250, -3660, -7402, 3358, 7537, -3057, -7659, 2754, 7766, -2454, -7861, 2154, 7941, -1858, -8011, 1563, 8067, -1273, -8113, 985, 8147, -704, -8172, 425, 8185, -153, -8191, -115, 8187, 376, -8176, -633, 8155, 882, -8130, -1126, 8095, 1362, -8057, -1593, 8011, 1816, -7962, -2034, 7906, 2243, -7848, -2447, 7785, 2642, -7720, -2832, 7651, 3014, -7581, -3190, 7507, 3358, -7434, -3522, 7357, 3676, -7282, -3826, 7204, 3968, -7127, -4105, 7049, 4234, -6974, -4359, 6897, 4476, -6823, -4589, 6748, 4694, -6677, -4795, 6605, 4889, -6538, -4980, 6470, 5063, -6407, -5143, 6344, 5216, -6286, -5287, 6229, 5350, -6176, -5410, 6125, 5464, -6079, -5516, 6034, 5561, -5995, -5603, 5957, 5639, -5924, -5674, 5893, 5701, -5868, -5727, 5845, 5747, -5828, -5765, 5812, 5777, -5802, -5786, 5794, 5790, -5793, -5792, 5793, 5788, -5798, -5782, 5806, 5771, -5820, -5757, 5835, 5737, -5857, -5715, 5880, 5687, -5909, -5657, 5940, 5621, -5976, -5583, 6013, 5538, -6057, -5491, 6101, 5437, -6151, -5381, 6202, 5318, -6258, -5253, 6314, 5180, -6376, -5104, 6438, 5022, -6504, -4936, 6571, 4842, -6641, -4746, 6712, 4641, -6786, -4533, 6859, 4417, -6936, -4298, 7011, 4170, -7089, -4038, 7165, 3897, -7243, -3752, 7319, 3599, -7396, -3441, 7470, 3275, -7545, -3103, 7616, 2923, -7687, -2738, 7753, 2544, -7818, -2346, 7877, 2138, -7935, -1926, 7987, 1705, -8035, -1479, 8076, 1244, -8114, -1005, 8143, 757, -8167, -505, 8182, 245, -8191, 18, 8189, -289, -8180, 564, 8160, -845, -8132, 1129, 8091, -1418, -8041, 1710, 7977, -2006, -7903, 2303, 7814, -2604, -7714, 2905, 7599, -3208, -7471, 3509, 7327, -3811, -7170, 4110, 6996, -4408, -6808, 4700, 6603, -4991, -6384, 5274, 6146, -5552, -5895, 5821, 5625, -6084, -5341, 6335, 5039, -6577, -4723, 6805, 4389, -7022, -4042, 7223, 3678, -7410, -3302, 7578, 2910, -7730, -2507, 7861, 2089, -7973, -1663, 8062, 1224, -8130, -778, 8172, 322, -8191, 138, 8182, -605, -8148, 1074, 8085, -1547, -7995, 2018, 7874, -2489, -7726, 2955, 7545, -3416, -7337, 3868, 7095, -4312, -6826, 4742, 6524, -5159, -6194, 5557, 5833, -5938, -5446, 6295, 5028, -6630, -4586, 6937, 4117, -7217, -3626, 7465, 3111, -7681, -2578, 7860, 2026, -8004, -1460, 8106, 879, -8171, -290, 8190, -309, -8169, 909, 8101, -1511, -7989, 2109, 7829, -2701, -7625, 3282, 7372, -3850, -7076, 4399, 6732, -4927, -6345, 5427, 5914, -5899, -5443, 6335, 4931, -6735, -4384, 7092, 3801, -7406, -3190, 7670, 2549, -7885, -1887, 8043, 1205, -8146, -510, 8189, -196, -8173, 904, 8093, -1612, -7953, 2312, 7747, -3001, -7481, 3669, 7150, -4314, -6761, 4927, 6311, -5506, -5806, 6040, 5246, -6528, -4639, 6960, 3985, -7337, -3292, 7648, 2563, -7894, -1807, 8067, 1027, -8167, -234, 8189, -569, -8134, 1369, 7997, -2164, -7783, 2941, 7487, -3695, -7115, 4415, 6665, -5095, -6145, 5725, 5554, -6300, -4902, 6808, 4191, -7248, -3431, 7608, 2626, -7888, -1788, 8077, 922, -8177, -42, 8181, -845, -8090, 1726, 7900, -2594, -7615, 3434, 7234, -4239, -6762, 4993, 6202, -5692, -5561, 6319, 4843, -6871, -4060, 7335, 3216, -7706, -2328, 7975, 1400, -8139, -450, 8190, -513, -8131, 1473, 7955, -2419, -7668, 3335, 7267, -4209, -6761, 5026, 6150, -5774, -5447, 6439, 4657, -7012, -3794, 7480, 2866, -7837, -1891, 8072, 878, -8183, 151, 8163, -1186, -8014, 2205, 7731, -3195, -7322, 4136, 6787, -5015, -6138, 5812, 5379, -6516, -4527, 7109, 3590, -7584, -2587, 7926, 1531, -8131, -445, 8190, -657, -8102, 1750, 7864, -2818, -7482, 3838, 6956, -4792, -6298, 5659, 5516, -6423, -4625, 7066, 3639, -7575, -2578, 7936, 1460, -8143, -309, 8186, -856, -8065, 2007, 7777, -3124, -7328, 4179, 6723, -5154, -5976, 6022, 5096, -6768, -4106, 7370, 3019, -7817, -1865, 8092, 661, -8191, 560, 8106, -1776, -7840, 2956, 7393, -4075, -6776, 5104, 5998, -6020, -5078, 6797, 4033, -7419, -2889, 7865, 1669, -8125, -406, 8187, -875, -8051, 2138, 7714, -3355, -7184, 4491, 6471, -5521, -5592, 6413, 4564, -7146, -3417, 7695, 2174, -8048, -871, 8188, -463, -8113, 1787, 7820, -3071, -7316, 4275, 6609, -5370, -5720, 6319, 4667, -7098, -3482, 7680, 2192, -8049, -837, 8189, -549, -8097, 1923, 7769, -3248, -7215, 4482, 6445, -5590, -5484, 6535, 4353, -7290, -3089, 7826, 1725, -8128, -304, 8180, -1132, -7982, 2538, 7533, -3871, -6847, 5086, 5941, -6146, -4845, 7012, 3587, -7657, -2211, 8054, 755, -8191, 729, 8058, -2196, -7659, 3593, 7000, -4877, -6105, 5999, 4999, -6923, -3719, 7611, 2305, -8041, -808, 8190, -725, -8056, 2235, 7634, -3674, -6942, 4985, 5997, -6124, -4834, 7043, 3490, -7710, -2015, 8096, 460, -8185, 1117, 7968, -2659, -7454, 4104, 6655, -5401, -5602, 6495, 4330, -7345, -2888, 7912, 1328, -8175, 288, 8116, -1900, -7740, 3440, 7053, -4850, -6083, 6068, 4863, -7047, -3445, 7741, 1879, -8122, -232, 8168, -1431, -7878, 3038, 7255, -4525, -6328, 5824, 5127, -6883, -3707, 7648, 2121, -8089, -441, 8180, -1266, -7917, 2921, 7303, -4455, -6368, 5795, 5144, -6882, -3689, 7663, 2062, -8102, -338, 8173, -1409, -7872, 3094, 7207, -4645, -6208, 5982, 4915, -7046, -3390, 7780, 1698, -8151, 77, 8133, -1856, -7727, 3550, 6946, -5079, -5828, 6363, 4421, -7343, -2794, 7962, 1023, -8191, 802, 8010, -2595, -7430, 4261, 6471, -5718, -5184, 6887, 3626, -7708, -1880, 8134, 29, -8141, 1827, 7723, -3594, -6901, 5176, 5711, -6491, -4216, 7462, 2491, -8039, -629, 8184, -1274, -7888, 3112, 7161, -4787, -6041, 6202, 4584, -7281, -2871, 7956, 991, -8191, 947, 7966, -2840, -7291, 4575, 6199, -6056, -4752, 7193, 3026, -7920, -1122, 8189, -854, -7984, 2783, 7309, -4557, -6203, 6064, 4725, -7217, -2964, 7941, 1019, -8191, 991, 7947, -2949, -7221, 4730, 6050, -6228, -4507, 7346, 2680, -8014, -684, 8183, -1362, -7844, 3326, 7008, -5087, -5729, 6529, 4081, -7561, -2170, 8109, 113, -8139, 1955, 7640, -3904, -6644, 5601, 5210, -6937, -3431, 7817, 1419, -8183, 691, 8003, -2762, -7289, 4651, 6081, -6232, -4460, 7393, 2529, -8055, -423, 8164, -1720, -7714, 3747, 6726, -5521, -5269, 6913, 3439, -7825, -1364, 8186, -815, -7970, 2939, 7184, -4860, -5884, 6436, 4156, -7553, -2125, 8124, -67, -8107, 2257, 7495, -4290, -6332, 6009, 4696, -7289, -2710, 8027, 514, -8169, 1723, 7695, -3838, -6640, 5665, 5077, -7068, -3125, 7931, 926, -8189, 1347, 7813, -3523, -6832, 5428, 5314, -6916, -3378, 7862, 1170, -8191, 1134, 7871, -3355, -6924, 5311, 5420, -6848, -3477, 7835, 1248, -8191, 1086, 7880, -3339, -6925, 5321, 5398, -6872, -3424, 7856, 1160, -8191, 1205, 7842, -3476, -6836, 5457, 5249, -6985, -3217, 7921, 905, -8186, 1488, 7749, -3761, -6647, 5712, 4965, -7175, -2851, 8015, 482, -8159, 1933, 7584, -4185, -6342, 6070, 4533, -7423, -2318, 8114, -110, -8082, 2532, 7321, -4733, -5898, 6508, 3935, -7696, -1610, 8182, -869, -7920, 3271, 6924, -5378, -5288, 6989, 3154, -7953, -723, 8173, -1783, -7627, 4125, 6357, -6083, -4484, 7465, 2177, -8139, 341, 8032, -2833, -7153, 5055, 5578, -6794, -3461, 7873, 999, -8187, 1564, 7695, -3980, -6445, 6006, 4553, -7442, -2206, 8137, -368, -8022, 2909, 7098, -5163, -5458, 6899, 3259, -7939, -726, 8169, -1888, -7566, 4312, 6181, -6298, -4157, 7635, 1695, -8183, 945, 7876, -3494, -6745, 5680, 4900, -7273, -2536, 8097, -104, -8064, 2736, 7169, -5083, -5505, 6886, 3243, -7953, -629, 8158, -2061, -7480, 4529, 5981, -6509, -3826, 7776, 1244, -8191, 1479, 7697, -4044, -6349, 6163, 4288, -7598, -1744, 8182, -1002, -7846, 3639, 6620, -5870, -4642, 7436, 2128, -8156, 632, 7941, -3327, -6812, 5641, 4891, -7308, -2401, 8126, -375, -7998, 3111, 6931, -5489, -5048, 7222, 2563, -8105, 228, 8025, -3000, -6990, 5416, 5113, -7189, -2620, 8097, -195, -8030, 2990, 6987, -5429, -5092, 7207, 2569, -8108, 272, 8011, -3087, -6927, 5523, 4980, -7280, -2412, 8130, -463, -7967, 3284, 6802, -5699, -4778, 7396, 2145, -8161, 764, 7887, -3583, -6607, 5946, 4476, -7552, -1767, 8185, -1177, -7762, 3972, 6329, -6257, -4070, 7727, 1273, -8189, 1695, 7572, -4446, -5957, 6612, 3547, -7906, -664, 8147, -2316, -7301, 4988, 5472, -6996, -2904, 8062, -63, -8040, 3025, 6922, -5581, -4861, 7378, 2129, -8168, 899, 7832, -3810, -6416, 6197, 4107, -7729, -1223, 8185, -1837, -7498, 4644, 5756, -6805, -3202, 8006, 189, -8078, 2854, 7000, -5498, -4924, 7359, 2138, -8169, 959, 7804, -3924, -6313, 6325, 3903, -7814, -924, 8165, -2198, -7325, 5000, 5408, -7075, -2693, 8108, -425, -7946, 3484, 6601, -6032, -4273, 7682, 1300, -8186, 1870, 7460, -4767, -5609, 6946, 2905, -8078, 243, 7982, -3360, -6670, 5968, 4332, -7666, -1328, 8186, -1889, -7444, 4816, 5546, -7003, -2785, 8101, -417, -7937, 3556, 6527, -6145, -4090, 7767, 1002, -8167, 2248, 7270, -5148, -5216, 7230, 2325, -8161, 941, 7782, -4064, -6152, 6534, 3524, -7953, -322, 8081, -2938, -6896, 5723, 4580, -7578, -1512, 8189, -1812, -7454, 4840, 5485, -7073, -2605, 8133, -715, -7842, 3919, 6238, -6473, -3587, 7943, 327, -8078, 2992, 6845, -5811, -4452, 7645, 1296, -8182, 2084, 7318, -5115, -5200, 7269, 2182, -8177, 1215, 7670, -4409, -5834, 6840, 2978, -8085, 400, 7916, -3715, -6361, 6380, 3682, -7927, -352, 8074, -3048, -6791, 5909, 4296, -7724, -1033, 8160, -2422, -7135, 5445, 4824, -7494, -1641, 8190, -1846, -7405, 5000, 5270, -7251, -2174, 8179, -1327, -7612, 4588, 5643, -7010, -2633, 8141, -871, -7767, 4215, 5948, -6783, -3020, 8086, -479, -7880, 3891, 6192, -6578, -3337, 8026, -154, -7960, 3619, 6382, -6403, -3588, 7969, 103, -8015, 3405, 6522, -6265, -3774, 7921, 292, -8050, 3249, 6618, -6167, -3898, 7886, 413, -8070, 3155, 6672, -6112, -3962, 7869, 467, -8077, 3124, 6686, -6103, -3967, 7870, 452, -8073, 3155, 6660, -6138, -3912, 7890, 370, -8057, 3249, 6595, -6218, -3796, 7927, 220, -8027, 3404, 6487, -6339, -3619, 7977, 2, -7978, 3618, 6333, -6498, -3378, 8035, -284, -7906, 3890, 6129, -6691, -3070, 8094, -637, -7803, 4214, 5868, -6910, -2694, 8147, -1057, -7661, 4586, 5545, -7146, -2245, 8182, -1540, -7471, 4999, 5152, -7389, -1723, 8188, -2084, -7220, 5443, 4683, -7627, -1127, 8151, -2682, -6899, 5908, 4132, -7844, -456, 8056, -3327, -6495, 6378, 3493, -8023, 285, 7887, -4007, -5997, 6838, 2763, -8146, 1092, 7627, -4709, -5395, 7268, 1941, -8191, 1954, 7260, -5413, -4681, 7644, 1031, -8137, 2857, 6769, -6098, -3850, 7942, 40, -7962, 3783, 6142, -6738, -2901, 8133, -1020, -7642, 4706, 5368, -7301, -1839, 8189, -2128, -7159, 5597, 4442, -7755, -676, 8082, -3257, -6497, 6421, 3365, -8064, 569, 7784, -4375, -5645, 7137, 2148, -8190, 1868, 7272, -5440, -4600, 7700, 809, -8100, 3180, 6530, -6403, -3370, 8066, -619, -7761, 4460, 5550, -7212, -1974, 8190, -2095, -7150, 5649, 4337, -7810, -447, 8031, -3562, -6254, 6685, 2911, -8142, 1164, 7557, -4953, -5074, 7498, 1307, -8155, 2793, 6748, -6192, -3629, 8021, -419, -7810, 4363, 5603, -7198, -1961, 8190, -2191, -7079, 5782, 4142, -7888, -132, 7953, -3918, -5958, 6954, 2410, -8185, 1769, 7279, -5493, -4469, 7780, 482, -8028, 3635, 6160, -6800, -2666, 8170, -1540, -7377, 5341, 4622, -7726, -634, 8052, -3530, -6227, 6752, 2729, -8167, 1505, 7384, -5340, -4611, 7736, 585, -8041, 3602, 6162, -6817, -2606, 8176, -1668, -7305, 5488, 4431, -7810, -338, 7986, -3854, -5963, 6985, 2289, -8190, 2021, 7124, -5777, -4078, 7928, -110, -7871, 4270, 5610, -7241, -1776, 8180, -2563, -6821, 6184, 3534, -8064, 755, 7660, -4836, -5084, 7545, 1056, -8110, 3275, 6358, -6677, -2785, 8167, -1593, -7314, 5515, 4351, -7854, -131, 7923, -4134, -5698, 7202, 1813, -8181, 2602, 6774, -6264, -3388, 8096, -997, -7557, 5091, 4793, -7694, -616, 8027, -3749, -5989, 7008, 2170, -8191, 2295, 6937, -6084, -3614, 8058, -794, -7624, 4968, 4900, -7656, -702, 8039, -3715, -5999, 7012, 2139, -8191, 2371, 6882, -6168, -3479, 8087, -990, -7541, 5160, 4683, -7755, -388, 7968, -4034, -5730, 7215, 1719, -8171, 2826, 6596, -6502, -2973, 8158, -1580, -7277, 5644, 4120, -7950, 327, 7765, -4679, -5142, 7562, 897, -8066, 3635, 6021, -7023, -2069, 8187, -2545, -6752, 6354, 3164, -8142, 1436, 7328, -5583, -4168, 7943, -335, -7754, 4733, 5065, -7611, -740, 8030, -3831, -5850, 7162, 1766, -8170, 2895, 6515, -6619, -2733, 8180, -1950, -7065, 5996, 3626, -8077, 1008, 7496, -5316, -4441, 7869, -90, -7818, 4593, 5169, -7576, -798, 8034, -3846, -5812, 7206, 1640, -8157, 3085, 6366, -6779, -2433, 8190, -2327, -6838, 6303, 3168, -8149, 1579, 7227, -5796, -3846, 8040, -853, -7542, 5263, 4460, -7876, 153, 7784, -4720, -5015, 7663, 511, -7965, 4172, 5508, -7416, -1140, 8086, -3630, -5945, 7139, 1727, -8160, 3098, 6325, -6844, -2273, 8189, -2585, -6656, 6535, 2773, -8184, 2092, 6938, -6223, -3232, 8147, -1626, -7178, 5909, 3647, -8089, 1188, 7377, -5604, -4022, 8012, -782, -7544, 5308, 4355, -7926, 407, 7679, -5029, -4652, 7830, -68, -7789, 4766, 4910, -7733, -238, 7876, -4527, -5136, 7636, 508, -7945, 4310, 5328, -7546, -745, 7997, -4120, -5491, 7461, 944, -8038, 3955, 5623, -7389, -1111, 8066, -3822, -5729, 7326, 1241, -8088, 3715, 5807, -7280, -1339, 8101, -3641, -5863, 7247, 1400, -8110, 3596, 5891, -7231, -1429, 8112, -3584, -5897, 7230, 1422, -8111, 3601, 5878, -7246, -1383, 8103, -3651, -5836, 7277, 1308, -8092, 3729, 5767, -7325, -1200, 8072, -3840, -5674, 7385, 1056, -8046, 3979, 5553, -7458, -879, 8008, -4147, -5405, 7541, 665, -7959, 4341, 5225, -7633, -418, 7894, -4562, -5016, 7728, 134, -7813, 4805, 4771, -7826, 183, 7708, -5071, -4493, 7920, -536, -7580, 5352, 4176, -8009, 921, 7421, -5650, -3821, 8085, -1340, -7231, 5957, 3423, -8146, 1787, 7001, -6270, -2985, 8182, -2263, -6730, 6582, 2501) 	  
    ) 
    port map (
    Clk_96 => Clk_96,
     Ce_F6 => Ce_F6,
     EN =>EN,
     Rom_cos_all => Rom_cos_L40C33_i
    );

process(Clk_96, Ce_F6 , TI , LG  )
    variable count: integer := 0;
    variable guard: boolean := False;
begin
    if TI = '1' then 	
	adress <= "11";
    elsif rising_edge(clk_96) then         
	    if LG = '0' and guard = False  then				 
		 guard := True;
		 adress <= adress +1;					 
		if adress = "11" then
		   adress <= "00";
		end if;
	    elsif LG = '1' then 
	       guard := False;
	    end if;	
    end if;					 
end process;

    pft_adress <= PFT & adress ;
process(PFT_adress, Rom_cos_L15_i, Rom_cos_L15�31_i, Rom_cos_L15�32_i, Rom_cos_L15�33_i, Rom_cos_L21_i, Rom_cos_L21C31_i, Rom_cos_L21C32_i, Rom_cos_L21C33_i, Rom_cos_L32_i, Rom_cos_L32C31_i, Rom_cos_L32C32_i, Rom_cos_L32C33_i, Rom_cos_L40_i, Rom_cos_L40C31_i, Rom_cos_L40C32_i, Rom_cos_L40C33_i)
begin
  if  pft_adress = "0110000000" or pft_adress = "0110001100" then
        Rom_cos_i <= Rom_cos_L15_i;
    elsif pft_adress = "0110000100" or pft_adress = "0110001000" or pft_adress = "0110011000" or pft_adress = "0110011100" or pft_adress = "0111000100" or pft_adress = "0111001000" or pft_adress = "0111011000" or pft_adress = "0111011100" then
        Rom_cos_i <= Rom_cos_L15�31_i;
    elsif pft_adress = "0110000101" or pft_adress = "0110001001" or pft_adress = "0110011001" or pft_adress = "0110011101" or pft_adress = "0111000101" or pft_adress = "0111001001" or pft_adress = "0111011001" or pft_adress = "0111011101" then
        Rom_cos_i <= Rom_cos_L15�32_i;
    elsif pft_adress = "0110000110" or pft_adress = "0110001010" or pft_adress = "0110011010" or pft_adress = "0110011110" or pft_adress = "0111000110" or pft_adress = "0111001010" or pft_adress = "0111011010" or pft_adress = "0111011110" then
        Rom_cos_i <= Rom_cos_L15�33_i;
    elsif pft_adress = "0100000000" or pft_adress = "0100001100" then
        Rom_cos_i <= Rom_cos_L21_i;
    elsif pft_adress = "0100000100" or pft_adress = "0100001000" or pft_adress = "0100011000" or pft_adress = "0100011100" or pft_adress = "0101000100" or pft_adress = "0101001000" or pft_adress = "0101011000" or pft_adress = "0101011100" then
        Rom_cos_i <= Rom_cos_L21C31_i;
    elsif pft_adress = "0100000101" or pft_adress = "0100001001" or pft_adress = "0100011001" or pft_adress = "0100011101" or pft_adress = "0101000101" or pft_adress = "0101001001" or pft_adress = "0101011001" or pft_adress = "0101011101" then
        Rom_cos_i <= Rom_cos_L21C32_i;
    elsif pft_adress = "0100000110" or pft_adress = "0100001010" or pft_adress = "0100011010" or pft_adress = "0100011110" or pft_adress = "0101000110" or pft_adress = "0101001010" or pft_adress = "0101011010" or pft_adress = "0101011110" then
        Rom_cos_i <= Rom_cos_L21C33_i;
    elsif pft_adress = "0010000000" or pft_adress = "0010001100" then
        Rom_cos_i <= Rom_cos_L32_i;
    elsif pft_adress = "0010000100" or pft_adress = "0010001000" or pft_adress = "0010011000" or pft_adress = "0010011100" or pft_adress = "0011000100" or pft_adress = "0011001000" or pft_adress = "0011011000" or pft_adress = "0011011100" then
        Rom_cos_i <= Rom_cos_L32C31_i;
    elsif pft_adress = "0010000101" or pft_adress = "0010001001" or pft_adress = "0010011001" or pft_adress = "0010011101" or pft_adress = "0011000101" or pft_adress = "0011001001" or pft_adress = "0011011001" or pft_adress = "0011011101" then
        Rom_cos_i <= Rom_cos_L32C32_i;
    elsif pft_adress = "0010000110" or pft_adress = "0010001010" or pft_adress = "0010011010" or pft_adress = "0010011110" or pft_adress = "0011000110" or pft_adress = "0011001010" or pft_adress = "0011011010" or pft_adress = "0011011110" then
        Rom_cos_i <= Rom_cos_L32C33_i;
    elsif pft_adress = "0000000000" or pft_adress = "0000001100" or pft_adress = "1100000000" then
        Rom_cos_i <= Rom_cos_L40_i;
    elsif pft_adress = "0000000100" or pft_adress = "0000001000" or pft_adress = "0000011000" or pft_adress = "0000011100" then
        Rom_cos_i <= Rom_cos_L40C31_i;
    elsif pft_adress = "0000000101" or pft_adress = "0000001001" or pft_adress = "0000011001" or pft_adress = "0000011101" then
        Rom_cos_i <= Rom_cos_L40C32_i;
    elsif pft_adress = "0000000110" or pft_adress = "0000001010" or pft_adress = "0000011010" or pft_adress = "0000011110" then
        Rom_cos_i <= Rom_cos_L40C33_i;
    end if; 
 end process;

process (Clk_96, Ce_F6, EN, Rom_cos_i )
begin
	 
    if EN = '1' then
       Rom_cos <= conv_std_logic_vector(Rom_cos_i- magic, data_rom);
    else
       Rom_cos <=(others => '0');
    end if;	
end process;end Behavioral;